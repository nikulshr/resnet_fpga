localparam BN12_CH = 64;
localparam BN12_BW_A = 6;
localparam BN12_BW_B = 15;
localparam BN12_RSHIFT = 8;
localparam BN12_BW_IN = 16;
localparam BN12_BW_OUT = 1;
localparam BN12_MAXVAL = 1;
reg [BN12_CH-1:0][BN12_BW_A-1:0] bn12_a = { 6'h10, 6'h11, 6'h0c, 6'h11, 6'h15, 6'h0c, 6'h19, 6'h0f, 6'h07, 6'h0e, 6'h18, 6'h10, 6'h0e, 6'h10, 6'h14, 6'h17, 6'h15, 6'h0f, 6'h13, 6'h15, 6'h0c, 6'h0f, 6'h0b, 6'h0b, 6'h16, 6'h13, 6'h13, 6'h11, 6'h14, 6'h13, 6'h10, 6'h14, 6'h17, 6'h17, 6'h13, 6'h12, 6'h0d, 6'h0c, 6'h14, 6'h0d, 6'h08, 6'h0d, 6'h0f, 6'h10, 6'h1f, 6'h15, 6'h09, 6'h0c, 6'h0c, 6'h1f, 6'h19, 6'h16, 6'h0e, 6'h17, 6'h0c, 6'h0f, 6'h0f, 6'h1c, 6'h11, 6'h15, 6'h12, 6'h09, 6'h11, 6'h13 };
reg [BN12_CH-1:0][BN12_BW_B-1:0] bn12_b = { 15'h1956, 15'h7823, 15'h01fb, 15'h16ae, 15'h68a5, 15'h7d80, 15'h16d2, 15'h782b, 15'h790d, 15'h14ce, 15'h1db8, 15'h7508, 15'h7d4b, 15'h1a0b, 15'h7ee7, 15'h6d16, 15'h1174, 15'h7ff1, 15'h5be1, 15'h6493, 15'h7aa1, 15'h7b0a, 15'h6f44, 15'h073c, 15'h17b2, 15'h66e7, 15'h1948, 15'h06ea, 15'h15ec, 15'h05f0, 15'h7004, 15'h13dd, 15'h7854, 15'h0b82, 15'h0144, 15'h7930, 15'h014d, 15'h60aa, 15'h087b, 15'h0000, 15'h6309, 15'h1124, 15'h1a72, 15'h0352, 15'h071f, 15'h7fde, 15'h6bfe, 15'h0582, 15'h0d3e, 15'h73ed, 15'h07d5, 15'h03c0, 15'h0acd, 15'h05e3, 15'h0327, 15'h0c12, 15'h0d23, 15'h063c, 15'h22fa, 15'h1a2b, 15'h089c, 15'h128f, 15'h15a8, 15'h0204 };
