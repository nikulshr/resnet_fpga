localparam D0_IN_SIZE = 2;
localparam D0_BW_W = 2;
localparam D0_SHIFT = 0;
localparam LOG2_D0_CYC = 6;
localparam D0_CYC = 64;
localparam D0_CH = 1024;
reg [LOG2_D0_CYC-1:0] d0_cntr;
wire [D0_CH-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0;
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_0 = { 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'hf, 4'h5, 4'hf, 4'h3, 4'hf, 4'h4, 4'hf, 4'h1, 4'hf, 4'h1, 4'h1, 4'h4, 4'hd, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'h1, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'hc, 4'h4, 4'h1, 4'h4, 4'h7, 4'h4, 4'h7, 4'hd, 4'hc, 4'hc, 4'h0, 4'h7, 4'h1, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'h7, 4'h0, 4'h3 };
assign dw_0[0] = dw_0_0[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1 = { 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h7, 4'h5, 4'h0, 4'hf, 4'hf, 4'h0, 4'hf, 4'h4, 4'hf, 4'hd, 4'hc, 4'h3, 4'h3, 4'h0, 4'h1, 4'hc, 4'hc, 4'h7, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'h3, 4'h4, 4'hc, 4'h0, 4'hc, 4'hf, 4'h3, 4'h4, 4'h1, 4'h0, 4'h4, 4'h3, 4'h3, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3 };
assign dw_0[1] = dw_0_1[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_2 = { 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h4, 4'hd, 4'h0, 4'h1, 4'h4, 4'h0, 4'hd, 4'h0, 4'h4, 4'hc, 4'h1, 4'h0, 4'hc, 4'h3, 4'h4, 4'hd, 4'h0, 4'h5, 4'hf, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h4 };
assign dw_0[2] = dw_0_2[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_3 = { 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h5, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'hc, 4'h0, 4'h4, 4'hd, 4'h0, 4'h1, 4'hf, 4'h3, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'hc, 4'hd, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3 };
assign dw_0[3] = dw_0_3[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_4 = { 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h7, 4'h5, 4'h0, 4'h0, 4'h3, 4'h4, 4'hf, 4'h7, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h7, 4'hc, 4'h4, 4'hc, 4'h4, 4'h0, 4'h3, 4'h4, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h1, 4'h5, 4'h1, 4'h0, 4'h1, 4'hf, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0 };
assign dw_0[4] = dw_0_4[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_5 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'h1, 4'h5, 4'h3, 4'h1, 4'h3, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd, 4'hc, 4'h4, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0 };
assign dw_0[5] = dw_0_5[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_6 = { 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h5, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'h4, 4'h3, 4'hc, 4'hf, 4'h0, 4'h3, 4'h5, 4'h1, 4'h0, 4'hc, 4'h7, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h1, 4'h4, 4'h3, 4'hd, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h5, 4'h3, 4'h3, 4'hd, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'hc, 4'h3, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0 };
assign dw_0[6] = dw_0_6[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_7 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h5, 4'h0, 4'h3, 4'hf, 4'h4, 4'hf, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h5, 4'hd, 4'h0, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0, 4'h4, 4'h3, 4'h5, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'h4, 4'h3, 4'hf, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0 };
assign dw_0[7] = dw_0_7[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_8 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h4, 4'h3, 4'hf, 4'h7, 4'hf, 4'h4, 4'hf, 4'h0, 4'hf, 4'h0, 4'h3, 4'h5, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h4, 4'h3, 4'h1, 4'hc, 4'hc, 4'h0, 4'h4, 4'hd, 4'h0, 4'h4, 4'hf, 4'h3, 4'h1, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0 };
assign dw_0[8] = dw_0_8[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_9 = { 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h7, 4'h5, 4'hc, 4'h0, 4'hf, 4'h4, 4'hf, 4'h4, 4'h3, 4'hc, 4'hc, 4'h3, 4'h3, 4'h4, 4'hd, 4'h0, 4'h0, 4'h3, 4'hc, 4'h4, 4'hc, 4'h5, 4'h0, 4'hf, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'h5, 4'h3, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h4, 4'h3, 4'h3, 4'h1, 4'hf, 4'h1, 4'h0, 4'h4, 4'hc, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'h4 };
assign dw_0[9] = dw_0_9[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_10 = { 4'h3, 4'h5, 4'h4, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h4, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h5, 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h5, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'hf, 4'h3, 4'hd, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0 };
assign dw_0[10] = dw_0_10[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_11 = { 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h7, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'hd, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0 };
assign dw_0[11] = dw_0_11[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_12 = { 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h3, 4'h4, 4'hf, 4'h3, 4'hf, 4'h7, 4'h3, 4'hd, 4'hf, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hd, 4'h0, 4'h3, 4'hc, 4'h5, 4'h1, 4'h0, 4'h5, 4'hf, 4'h3, 4'h1, 4'hf, 4'h7, 4'h0, 4'h3, 4'hc, 4'hf, 4'hd, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0 };
assign dw_0[12] = dw_0_12[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_13 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'h5, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'h4, 4'h3, 4'hc, 4'hc, 4'h3, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'hf, 4'h1, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'h3, 4'h3, 4'hd, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0 };
assign dw_0[13] = dw_0_13[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_14 = { 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h1, 4'h3, 4'hf, 4'h3, 4'hf, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h1, 4'hc, 4'h0, 4'h4, 4'hc, 4'hd, 4'hc, 4'h1, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'hf, 4'h3, 4'h1, 4'hf, 4'h0, 4'h0, 4'h7, 4'hc, 4'hf, 4'h1, 4'hc, 4'h0, 4'h0, 4'h1, 4'hf, 4'h4, 4'h4 };
assign dw_0[14] = dw_0_14[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_15 = { 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h5, 4'hf, 4'hc, 4'hf, 4'h7, 4'hc, 4'hc, 4'hc, 4'h1, 4'h1, 4'h3, 4'h1, 4'h0, 4'h4, 4'hf, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h4, 4'h4, 4'hd, 4'h0, 4'hc, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hd, 4'hd, 4'hc, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0 };
assign dw_0[15] = dw_0_15[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_16 = { 4'h5, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'h3, 4'hc, 4'h3, 4'h0, 4'hc, 4'h5, 4'h0, 4'hd, 4'h3, 4'h4, 4'h3, 4'h3, 4'h3, 4'h0, 4'hd, 4'h0, 4'h1, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h4, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc };
assign dw_0[16] = dw_0_16[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_17 = { 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'hc, 4'h5, 4'h0, 4'hd, 4'h3, 4'h0, 4'h7, 4'h1, 4'h0, 4'h3, 4'h1, 4'hc, 4'hd, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h0, 4'hc, 4'hd, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'hc, 4'h4, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h3, 4'h3, 4'h0, 4'h1, 4'h1, 4'h0, 4'hf };
assign dw_0[17] = dw_0_17[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_18 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'h1, 4'h1, 4'h5, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h7, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf };
assign dw_0[18] = dw_0_18[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_19 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hd, 4'hd, 4'hc, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h4, 4'h3, 4'h3, 4'hf, 4'h4, 4'h0, 4'hc, 4'h1, 4'h1, 4'h3, 4'h4, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'h4, 4'hc };
assign dw_0[19] = dw_0_19[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_20 = { 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h5, 4'h3, 4'h5, 4'h0, 4'hc, 4'h7, 4'hf, 4'h4, 4'h0, 4'hc, 4'h3, 4'hd, 4'hc, 4'hd, 4'hc, 4'h3, 4'h3, 4'h1, 4'h0, 4'h1, 4'h7, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h4, 4'h3, 4'h4, 4'h7, 4'h0, 4'hf, 4'h7, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'h0, 4'hc };
assign dw_0[20] = dw_0_20[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_21 = { 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h4, 4'h0, 4'h5, 4'h0, 4'h1, 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'hd, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'hd, 4'h3, 4'h3, 4'hc, 4'hf, 4'h3, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'h4, 4'h4, 4'h3, 4'hf, 4'h7, 4'h0, 4'h1, 4'h1, 4'h1, 4'hf, 4'h4, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hd, 4'h0, 4'h4, 4'hc };
assign dw_0[21] = dw_0_21[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_22 = { 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h5, 4'h0, 4'h5, 4'h4, 4'hd, 4'h4, 4'h3, 4'h3, 4'h3, 4'h7, 4'h3, 4'h0, 4'hc, 4'hd, 4'hc, 4'h3, 4'h3, 4'h1, 4'h0, 4'hc, 4'h3, 4'h7, 4'h3, 4'hf, 4'hf, 4'h0, 4'hc, 4'h1, 4'hf, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0, 4'hc, 4'h1, 4'h1, 4'hf, 4'h4, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc };
assign dw_0[22] = dw_0_22[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_23 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h5, 4'h3, 4'h5, 4'h0, 4'hc, 4'h3, 4'hc, 4'h4, 4'h3, 4'hf, 4'h3, 4'h0, 4'hc, 4'h1, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'hd, 4'h3, 4'h5, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc };
assign dw_0[23] = dw_0_23[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_24 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'hc, 4'h5, 4'h0, 4'hd, 4'h7, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'hc, 4'hd, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'hd, 4'h7, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'h0, 4'hc, 4'h7, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hf, 4'h7, 4'h0, 4'hc, 4'h5, 4'h4, 4'hf, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'hf };
assign dw_0[24] = dw_0_24[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_25 = { 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'hc, 4'h5, 4'h0, 4'hd, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'hc, 4'hd, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'hf, 4'h7, 4'h0, 4'h0, 4'h5, 4'h1, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'hc };
assign dw_0[25] = dw_0_25[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_26 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'hd, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h5, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'hf, 4'h7, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf };
assign dw_0[26] = dw_0_26[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_27 = { 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'hf, 4'h3, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h7, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc };
assign dw_0[27] = dw_0_27[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_28 = { 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hd, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'hc, 4'hc, 4'hc, 4'h0, 4'hc, 4'hf, 4'hc, 4'h0, 4'h4, 4'h4, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'hf };
assign dw_0[28] = dw_0_28[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_29 = { 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h7, 4'hc, 4'h0, 4'h3, 4'h5, 4'h0, 4'h5, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'hc };
assign dw_0[29] = dw_0_29[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_30 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h5, 4'h0, 4'hc, 4'h7, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'hc, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h7, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'hf, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h4, 4'hc };
assign dw_0[30] = dw_0_30[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_31 = { 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'hc, 4'hd, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h1, 4'hc, 4'hf, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h3, 4'hd, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h7, 4'h0, 4'hf, 4'h1, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf };
assign dw_0[31] = dw_0_31[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_32 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'hd, 4'h3, 4'h0, 4'h3, 4'h1, 4'h3, 4'h1, 4'hc, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h7, 4'hd, 4'h1, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0, 4'h7, 4'hc, 4'hf, 4'hc, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[32] = dw_0_32[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_33 = { 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h3, 4'h1, 4'hc, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h5, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'hf, 4'hc, 4'hf, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'hc, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0 };
assign dw_0[33] = dw_0_33[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_34 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h5, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h7, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0 };
assign dw_0[34] = dw_0_34[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_35 = { 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'h1, 4'h0, 4'h0, 4'hd, 4'h3, 4'h5, 4'h3, 4'hc, 4'h3, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'hc, 4'h0, 4'hd, 4'hf, 4'h0, 4'hf, 4'hd, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h7, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[35] = dw_0_35[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_36 = { 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc, 4'h5, 4'h0, 4'h4, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'h3, 4'h4, 4'h3, 4'h7, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'hd, 4'h5, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'hf, 4'hc, 4'hf, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'h5, 4'h7, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0 };
assign dw_0[36] = dw_0_36[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_37 = { 4'h1, 4'h5, 4'hc, 4'h1, 4'h0, 4'h4, 4'hc, 4'h1, 4'h4, 4'h4, 4'h1, 4'h3, 4'h4, 4'h3, 4'hd, 4'hf, 4'h5, 4'h3, 4'h4, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h1, 4'h3, 4'hd, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'hc, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h4, 4'h0 };
assign dw_0[37] = dw_0_37[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_38 = { 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h1, 4'h0, 4'h4, 4'hc, 4'h0, 4'h5, 4'h0, 4'hd, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'h5, 4'hc, 4'h3, 4'h0, 4'hd, 4'h1, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'hc, 4'h3, 4'hd, 4'h4, 4'h4, 4'h1, 4'h1, 4'h0, 4'hd, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0 };
assign dw_0[38] = dw_0_38[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_39 = { 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc, 4'h1, 4'hc, 4'h0, 4'h0, 4'h7, 4'h5, 4'h3, 4'h1, 4'hf, 4'h7, 4'h3, 4'h3, 4'h0, 4'h5, 4'hc, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0 };
assign dw_0[39] = dw_0_39[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_40 = { 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc, 4'h7, 4'h4, 4'h3, 4'h1, 4'hf, 4'h7, 4'h3, 4'h0, 4'h0, 4'h1, 4'hd, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'hd, 4'hc, 4'hc, 4'hf, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hd, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h5, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[40] = dw_0_40[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_41 = { 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h3, 4'h1, 4'hf, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'hc, 4'h3, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc, 4'h3, 4'hc, 4'hf, 4'hd, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h1, 4'hc, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h7, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0 };
assign dw_0[41] = dw_0_41[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_42 = { 4'h5, 4'h5, 4'h0, 4'h3, 4'h0, 4'h4, 4'hf, 4'hd, 4'h0, 4'h7, 4'h1, 4'h3, 4'h5, 4'h3, 4'h1, 4'hf, 4'h4, 4'h3, 4'h7, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'hd, 4'h1, 4'h4, 4'h0, 4'hc, 4'h4, 4'h7, 4'h7, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'h4, 4'h0, 4'h0, 4'h7, 4'h7, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h1, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h4 };
assign dw_0[42] = dw_0_42[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_43 = { 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h4, 4'hf, 4'hc, 4'hf, 4'h7, 4'h3, 4'h5, 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'h1, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'h3, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h4, 4'h0 };
assign dw_0[43] = dw_0_43[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_44 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'hd, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'hc, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'hd, 4'h4, 4'h0, 4'h1, 4'hc, 4'hc, 4'hc, 4'hc, 4'hc, 4'hf, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0 };
assign dw_0[44] = dw_0_44[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_45 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'h1, 4'h0, 4'hc, 4'h0, 4'h4, 4'hf, 4'hc, 4'h3, 4'h1, 4'h0, 4'h7, 4'h1, 4'h0, 4'hc, 4'h3, 4'hc, 4'hc, 4'h3, 4'h4, 4'h0, 4'h1, 4'h4, 4'h4, 4'h4, 4'hd, 4'h1, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'hf, 4'hc, 4'hf, 4'hd, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hf, 4'h5, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0 };
assign dw_0[45] = dw_0_45[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_46 = { 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'hd, 4'h3, 4'h0, 4'h0, 4'h7, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hd, 4'hd, 4'hc, 4'h0, 4'hf, 4'hc, 4'hf, 4'hd, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h5, 4'h7, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc };
assign dw_0[46] = dw_0_46[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_47 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'hc, 4'h1, 4'hf, 4'hc, 4'hf, 4'hc, 4'hd, 4'h7, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0 };
assign dw_0[47] = dw_0_47[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_48 = { 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h5, 4'h4, 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'hc, 4'h5, 4'h4, 4'hf, 4'h0, 4'hc, 4'hd, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h7, 4'h0, 4'h1, 4'h7, 4'hf, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'hf, 4'hc, 4'h4, 4'h0, 4'h5, 4'hf, 4'h4, 4'h1, 4'h3, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h5 };
assign dw_0[48] = dw_0_48[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_49 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3, 4'h7, 4'h0, 4'h7, 4'h0, 4'hd, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h1, 4'h5, 4'h4, 4'hd, 4'h3, 4'hc, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h7, 4'h0, 4'h3, 4'h7, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h5, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4 };
assign dw_0[49] = dw_0_49[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_50 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'hd, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h5, 4'h5, 4'hc, 4'h3, 4'hd, 4'hc, 4'hc, 4'hc, 4'h7, 4'hc, 4'hf, 4'hc, 4'h0, 4'h7, 4'h0, 4'h7, 4'h7, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'hc, 4'h0 };
assign dw_0[50] = dw_0_50[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_51 = { 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h1, 4'h4, 4'h5, 4'hd, 4'h3, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'hf, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1 };
assign dw_0[51] = dw_0_51[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_52 = { 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'hd, 4'h3, 4'h1, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'hd, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h4, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h1, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'hc, 4'h4 };
assign dw_0[52] = dw_0_52[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_53 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hd, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd, 4'h0, 4'h5, 4'h5, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'hc, 4'hf, 4'hd, 4'h1, 4'h3, 4'h0, 4'h3, 4'h7, 4'h3, 4'h0, 4'hd, 4'h4, 4'h0, 4'h1, 4'h3, 4'h7, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0 };
assign dw_0[53] = dw_0_53[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_54 = { 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'hd, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'hd, 4'h4, 4'h5, 4'hd, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'h3, 4'hc, 4'hf, 4'hd, 4'h5, 4'h7, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h1, 4'h3, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'hc, 4'h0 };
assign dw_0[54] = dw_0_54[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_55 = { 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h1, 4'h5, 4'h5, 4'hc, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5 };
assign dw_0[55] = dw_0_55[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_56 = { 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hd, 4'h4, 4'h4, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'h7, 4'h3, 4'h4, 4'hc, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'hc, 4'h5 };
assign dw_0[56] = dw_0_56[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_57 = { 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h1, 4'h3, 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h7, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'h1, 4'h4, 4'h1, 4'h3, 4'h7, 4'h0, 4'h4, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4 };
assign dw_0[57] = dw_0_57[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_58 = { 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h1, 4'h5, 4'h5, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h5 };
assign dw_0[58] = dw_0_58[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_59 = { 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'h1, 4'h4, 4'h5, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h4, 4'h0, 4'h1, 4'h3, 4'h7, 4'h3, 4'h5, 4'h1, 4'h7, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h4 };
assign dw_0[59] = dw_0_59[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_60 = { 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd, 4'h3, 4'h3, 4'h1, 4'h4, 4'h0, 4'h3, 4'h1, 4'h3, 4'hd, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd, 4'hd, 4'h5, 4'h5, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h3, 4'hc, 4'hf, 4'h1, 4'h0, 4'h7, 4'h0, 4'h7, 4'h4, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'hc, 4'h4 };
assign dw_0[60] = dw_0_60[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_61 = { 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'hd, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h7, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h4, 4'hc, 4'h3, 4'h1, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'hf, 4'hc, 4'h4, 4'h4, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h7, 4'h4, 4'h1, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'hd, 4'h0, 4'h1 };
assign dw_0[61] = dw_0_61[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_62 = { 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'hc, 4'h3, 4'h1, 4'h0, 4'h1, 4'h3, 4'hd, 4'h0, 4'h3, 4'h3, 4'hc, 4'hc, 4'h4, 4'h0, 4'h3, 4'h4, 4'hd, 4'h1, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'h4, 4'hc, 4'h3, 4'hc, 4'h0, 4'h1, 4'hc, 4'h7, 4'hc, 4'hf, 4'h1, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h5, 4'hc, 4'h4, 4'h0, 4'h1, 4'h7, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4 };
assign dw_0[62] = dw_0_62[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_63 = { 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h5, 4'hc, 4'h1, 4'hc, 4'h4, 4'h1, 4'hf, 4'h4, 4'h3, 4'h1, 4'h0, 4'h7, 4'h3, 4'h3, 4'h3, 4'h7, 4'h1, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hd, 4'h4, 4'h4, 4'hd, 4'h3, 4'hc, 4'hc, 4'h1, 4'hf, 4'h4, 4'hc, 4'hf, 4'hd, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h7, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h7, 4'h3, 4'hc, 4'h0 };
assign dw_0[63] = dw_0_63[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_64 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'h4, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h7, 4'h7, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'h0, 4'h7, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0 };
assign dw_0[64] = dw_0_64[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_65 = { 4'h0, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h4, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h4, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h7, 4'h3, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc };
assign dw_0[65] = dw_0_65[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_66 = { 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'h3, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h1, 4'h4, 4'h3, 4'h0, 4'h7, 4'h3, 4'h0, 4'h1, 4'h3, 4'hd, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0 };
assign dw_0[66] = dw_0_66[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_67 = { 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'hd, 4'hf, 4'hc, 4'h0, 4'hd, 4'h3, 4'h4, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h1, 4'h4, 4'h4, 4'hd, 4'h0, 4'hf, 4'h5, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'hd, 4'h3, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0 };
assign dw_0[67] = dw_0_67[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_68 = { 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'hd, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h4, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h1, 4'h7, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0 };
assign dw_0[68] = dw_0_68[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_69 = { 4'h0, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'hf, 4'h4, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'h1, 4'h0, 4'h3, 4'h0, 4'h7, 4'h3, 4'h0, 4'h1, 4'h1, 4'hd, 4'h0, 4'h0, 4'hf, 4'h7, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0 };
assign dw_0[69] = dw_0_69[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_70 = { 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'hf, 4'h5, 4'h0, 4'h3, 4'hf, 4'hc, 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'h7, 4'h7, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[70] = dw_0_70[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_71 = { 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h7, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h1, 4'h1, 4'h0, 4'hd, 4'h0, 4'h1, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0 };
assign dw_0[71] = dw_0_71[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_72 = { 4'h0, 4'hc, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h4, 4'h0, 4'h0, 4'hd, 4'h3, 4'hf, 4'h5, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h7, 4'h3, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1 };
assign dw_0[72] = dw_0_72[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_73 = { 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'hf, 4'hc, 4'h1, 4'h0, 4'h7, 4'h0, 4'hf, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'hf, 4'h1, 4'h0, 4'h0, 4'hd, 4'h0, 4'hf, 4'h5, 4'h4, 4'h3, 4'hc, 4'hc, 4'hc, 4'h3, 4'h4, 4'h3, 4'h0, 4'h7, 4'h3, 4'h1, 4'h5, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[73] = dw_0_73[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_74 = { 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'hf, 4'h1, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h7, 4'h7, 4'h0, 4'h5, 4'h0, 4'hd, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0 };
assign dw_0[74] = dw_0_74[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_75 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h1, 4'h5, 4'hd, 4'h0, 4'hf, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'h0, 4'h3, 4'h4, 4'h0, 4'h5, 4'h0, 4'hd, 4'h0, 4'h1, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc };
assign dw_0[75] = dw_0_75[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_76 = { 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'hd, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h1, 4'h3, 4'hc, 4'h1, 4'h3, 4'hc, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hd, 4'h3, 4'hf, 4'h4, 4'hf, 4'h3, 4'h3, 4'hc, 4'h3, 4'hc, 4'h4, 4'h3, 4'h0, 4'h7, 4'h4, 4'h0, 4'h5, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h7, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1 };
assign dw_0[76] = dw_0_76[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_77 = { 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'hd, 4'h0, 4'hf, 4'h5, 4'h3, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h7, 4'h7, 4'h0, 4'h5, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[77] = dw_0_77[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_78 = { 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h0, 4'h4, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h4, 4'hd, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h7, 4'h4, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'h7, 4'h5, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0 };
assign dw_0[78] = dw_0_78[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_79 = { 4'h3, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'hd, 4'h0, 4'h3, 4'h4, 4'hf, 4'h7, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc };
assign dw_0[79] = dw_0_79[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_80 = { 4'h0, 4'hf, 4'h4, 4'h3, 4'h0, 4'hc, 4'hf, 4'h3, 4'h5, 4'h1, 4'h1, 4'h5, 4'h0, 4'hd, 4'h7, 4'h0, 4'hf, 4'h1, 4'hd, 4'h1, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'hc, 4'h4, 4'h1, 4'hc, 4'hf, 4'hc, 4'h3, 4'hc, 4'h3, 4'h7, 4'h1, 4'h7, 4'hc, 4'hf, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h7, 4'h1, 4'h0, 4'hc, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h1, 4'hc, 4'hc };
assign dw_0[80] = dw_0_80[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_81 = { 4'h0, 4'hf, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h1, 4'h1, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hd, 4'h1, 4'h3, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'h3, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h7, 4'h1, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0 };
assign dw_0[81] = dw_0_81[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_82 = { 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'hd, 4'h1, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h3, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hd, 4'hf, 4'h1, 4'h3, 4'hc, 4'h3, 4'hf, 4'h5, 4'h4, 4'h3, 4'h7, 4'h4, 4'h3, 4'h1, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'h3, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0 };
assign dw_0[82] = dw_0_82[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_83 = { 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'hc, 4'hd, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'h1, 4'h7, 4'h0, 4'h4, 4'h4, 4'h4, 4'h5, 4'hc, 4'hf, 4'h0, 4'h7, 4'h0, 4'h0, 4'hd, 4'h4, 4'hc, 4'h0, 4'h0, 4'h7, 4'h4, 4'h5, 4'h7, 4'h0, 4'h0, 4'h5, 4'h3, 4'hc, 4'h0 };
assign dw_0[83] = dw_0_83[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_84 = { 4'h3, 4'hc, 4'h4, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h0, 4'hc, 4'h3, 4'hf, 4'h3, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'hd, 4'h7, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'hf, 4'h0, 4'h3, 4'h1, 4'hd, 4'hd, 4'h5, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h7, 4'h1, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc };
assign dw_0[84] = dw_0_84[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_85 = { 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'hd, 4'h0, 4'h3, 4'hc, 4'h5, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'h5, 4'h4, 4'h0, 4'h4, 4'h4, 4'h7, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h4, 4'h3, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[85] = dw_0_85[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_86 = { 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h1, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'hd, 4'h3, 4'h3, 4'h0, 4'h5, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'hc, 4'h1, 4'h7, 4'h0, 4'h7, 4'h4, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h7, 4'h1, 4'h0, 4'h5, 4'h4, 4'h3, 4'h0, 4'h0, 4'h7, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'hc };
assign dw_0[86] = dw_0_86[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_87 = { 4'h3, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h1, 4'h0, 4'hd, 4'h3, 4'h3, 4'h0, 4'h1, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'hc, 4'h7, 4'hf, 4'h3, 4'h3, 4'h1, 4'h7, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h7, 4'hc, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'h7, 4'hc, 4'h7, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0 };
assign dw_0[87] = dw_0_87[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_88 = { 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hd, 4'h1, 4'h5, 4'h7, 4'h1, 4'h3, 4'h3, 4'h1, 4'h3, 4'hd, 4'h1, 4'hf, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'hc, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h7, 4'h3, 4'h1, 4'h4, 4'h4, 4'h3, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4, 4'h5, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0 };
assign dw_0[88] = dw_0_88[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_89 = { 4'h3, 4'hc, 4'h4, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h4, 4'h0, 4'h3, 4'h3, 4'h1, 4'h3, 4'hd, 4'h1, 4'h3, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h7, 4'h0, 4'h4, 4'h4, 4'h3, 4'h7, 4'h3, 4'h3, 4'h0, 4'h7, 4'h0, 4'h3, 4'h4, 4'h5, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'hc, 4'h0 };
assign dw_0[89] = dw_0_89[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_90 = { 4'h3, 4'hd, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'hd, 4'h3, 4'h3, 4'h1, 4'h3, 4'h1, 4'h0, 4'h3, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'hd, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h7, 4'h4, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h7, 4'h1, 4'h0, 4'h4, 4'h5, 4'hf, 4'h0, 4'h0, 4'h7, 4'h4, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0 };
assign dw_0[90] = dw_0_90[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_91 = { 4'h3, 4'hc, 4'h4, 4'h3, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'hd, 4'h4, 4'h0, 4'hc, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h7, 4'h3, 4'h0, 4'h0, 4'h1, 4'hd, 4'hf, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[91] = dw_0_91[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_92 = { 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'h1, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'h3, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hd, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'h4, 4'h7, 4'h0, 4'h3, 4'h4, 4'h5, 4'h1, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h3, 4'h4, 4'h4, 4'hf, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'hc };
assign dw_0[92] = dw_0_92[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_93 = { 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'hd, 4'h3, 4'h0, 4'h5, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'h1, 4'hd, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h5, 4'h7, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h7, 4'h1, 4'h3, 4'h4, 4'h4, 4'hf, 4'h0, 4'h0, 4'h7, 4'h4, 4'hc, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0 };
assign dw_0[93] = dw_0_93[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_94 = { 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'hd, 4'h1, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h5, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'h3, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h5, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h7, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0 };
assign dw_0[94] = dw_0_94[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_95 = { 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'hd, 4'h0, 4'hf, 4'h0, 4'h5, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'hc, 4'h3, 4'hf, 4'h3, 4'h3, 4'h5, 4'h7, 4'h0, 4'h3, 4'h4, 4'h4, 4'h5, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[95] = dw_0_95[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_96 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h4, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h5, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'h7, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h5, 4'h0, 4'h1, 4'hc, 4'h5, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[96] = dw_0_96[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_97 = { 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'h1, 4'h1, 4'h3, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'h7, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h5, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h3, 4'h0, 4'h4, 4'hf, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'hc, 4'h4, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h3 };
assign dw_0[97] = dw_0_97[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_98 = { 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'h1, 4'hf, 4'h3, 4'h3, 4'h3, 4'h3, 4'h0, 4'hd, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h3, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hf, 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'hc, 4'h5, 4'h0, 4'h1, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0 };
assign dw_0[98] = dw_0_98[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_99 = { 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'hd, 4'h1, 4'hf, 4'h3, 4'h3, 4'hf, 4'hc, 4'hd, 4'hc, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[99] = dw_0_99[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_100 = { 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'hc, 4'h0, 4'hc, 4'hc, 4'h1, 4'h1, 4'h3, 4'h3, 4'h3, 4'hc, 4'h3, 4'h1, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'hd, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'hc, 4'h4, 4'h1, 4'h4, 4'h5, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0 };
assign dw_0[100] = dw_0_100[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_101 = { 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h1, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'hd, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h1, 4'hc, 4'h7, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[101] = dw_0_101[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_102 = { 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'hd, 4'h1, 4'h1, 4'h3, 4'h7, 4'h0, 4'h3, 4'h0, 4'h1, 4'hd, 4'h7, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'hc, 4'h4, 4'hf, 4'h1, 4'hc, 4'h7, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[102] = dw_0_102[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_103 = { 4'h4, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'h1, 4'h1, 4'h0, 4'hd, 4'hd, 4'h1, 4'hf, 4'h7, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h7, 4'hd, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'hf, 4'h1, 4'hc, 4'h4, 4'h0, 4'h3, 4'h5, 4'h4, 4'h0, 4'hc, 4'h5, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h3, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0 };
assign dw_0[103] = dw_0_103[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_104 = { 4'h4, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'hc, 4'hd, 4'h1, 4'h1, 4'hf, 4'h7, 4'h3, 4'hf, 4'h0, 4'h0, 4'hd, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'hd, 4'h3, 4'h5, 4'h1, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'h1, 4'hc, 4'h7, 4'h1, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h7, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[104] = dw_0_104[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_105 = { 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'h1, 4'h0, 4'h0, 4'hd, 4'h1, 4'h1, 4'h3, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'hc, 4'h7, 4'h1, 4'h0, 4'h5, 4'h1, 4'h3, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[105] = dw_0_105[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_106 = { 4'h4, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'hc, 4'hd, 4'h1, 4'h5, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'h5, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0 };
assign dw_0[106] = dw_0_106[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_107 = { 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h1, 4'h0, 4'hc, 4'hd, 4'h1, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'h7, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'hd, 4'h3, 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h1, 4'hc, 4'h7, 4'h0, 4'h0, 4'h5, 4'h4, 4'hc, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0 };
assign dw_0[107] = dw_0_107[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_108 = { 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'h1, 4'h3, 4'h3, 4'h0, 4'h3, 4'h3, 4'h1, 4'hc, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0 };
assign dw_0[108] = dw_0_108[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_109 = { 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h1, 4'hd, 4'hc, 4'h1, 4'h1, 4'h3, 4'h7, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h4, 4'hf, 4'h1, 4'hc, 4'h7, 4'h0, 4'h3, 4'h5, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h3, 4'h0, 4'hd, 4'h3, 4'h5, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0 };
assign dw_0[109] = dw_0_109[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_110 = { 4'h4, 4'hd, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'h1, 4'h3, 4'h0, 4'hd, 4'h0, 4'hc, 4'hd, 4'h5, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h1, 4'hc, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'hf, 4'h1, 4'hc, 4'h7, 4'h0, 4'h7, 4'h5, 4'h0, 4'hc, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h5, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[110] = dw_0_110[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_111 = { 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'hc, 4'hd, 4'h0, 4'hc, 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'h1, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h1, 4'h1, 4'h4, 4'h1, 4'h0, 4'h5, 4'h4, 4'hc, 4'hc, 4'h4, 4'h0, 4'h1, 4'h3, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0 };
assign dw_0[111] = dw_0_111[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_112 = { 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h7, 4'hc, 4'hf, 4'h4, 4'h4, 4'h3, 4'h1, 4'h1, 4'h0, 4'h5, 4'h4, 4'h0, 4'hd, 4'hc, 4'h3, 4'hc, 4'h0, 4'h4, 4'h4, 4'h4, 4'h3, 4'h1, 4'hd, 4'h4, 4'hc, 4'h7, 4'hf, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'h1, 4'hc, 4'h1, 4'h3, 4'hf, 4'hd, 4'h3, 4'hf, 4'h0, 4'h5, 4'h0, 4'h7, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'hf, 4'h4, 4'h5 };
assign dw_0[112] = dw_0_112[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_113 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hd, 4'hc, 4'h7, 4'h3, 4'hf, 4'h0, 4'hd, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h4, 4'h0, 4'h5, 4'h7, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h1, 4'h5, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hc, 4'h5, 4'hc, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h3, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hd, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc };
assign dw_0[113] = dw_0_113[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_114 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'hf, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h4, 4'h5, 4'h3, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'hc, 4'hf, 4'h0, 4'h3, 4'hc, 4'hc, 4'hf, 4'hd, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h7, 4'h0, 4'hc, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0 };
assign dw_0[114] = dw_0_114[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_115 = { 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h5, 4'h4, 4'h5, 4'h3, 4'h4, 4'h3, 4'hf, 4'h0, 4'h4, 4'hc, 4'h1, 4'h4, 4'hc, 4'hc, 4'h7, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h7, 4'h3, 4'h1, 4'h0, 4'h4, 4'h3, 4'h4, 4'h3 };
assign dw_0[115] = dw_0_115[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_116 = { 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'h7, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'h1, 4'h0, 4'hf, 4'h5, 4'h4, 4'h5, 4'h3, 4'h4, 4'hf, 4'hc, 4'hc, 4'h0, 4'hc, 4'h1, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'hc, 4'hc, 4'h1, 4'h1, 4'hc, 4'h4, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'hf, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'h7, 4'h3, 4'hc, 4'hf };
assign dw_0[116] = dw_0_116[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_117 = { 4'h3, 4'hd, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h3, 4'h0, 4'h5, 4'h4, 4'h5, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h4, 4'h0, 4'hc, 4'h4, 4'h0, 4'hc, 4'h1, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0 };
assign dw_0[117] = dw_0_117[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_118 = { 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'h7, 4'h0, 4'hf, 4'h4, 4'h0, 4'hc, 4'h3, 4'h1, 4'h0, 4'hc, 4'h5, 4'h4, 4'h5, 4'h4, 4'h4, 4'h3, 4'hc, 4'hc, 4'h0, 4'hc, 4'hc, 4'h5, 4'h0, 4'hc, 4'h4, 4'h3, 4'hc, 4'hc, 4'hf, 4'h0, 4'h4, 4'hc, 4'hd, 4'h1, 4'hc, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'h0, 4'h0 };
assign dw_0[118] = dw_0_118[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_119 = { 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'hc, 4'h1, 4'h7, 4'h0, 4'hf, 4'h5, 4'h1, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h4, 4'h0, 4'h5, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0 };
assign dw_0[119] = dw_0_119[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_120 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h5, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'hd, 4'hc, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'h0, 4'h0 };
assign dw_0[120] = dw_0_120[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_121 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'hf, 4'h4, 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'hc, 4'h1, 4'h4, 4'h4, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h1, 4'hc, 4'h1, 4'h1, 4'h3, 4'h7, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3 };
assign dw_0[121] = dw_0_121[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_122 = { 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'h3, 4'h4, 4'hc, 4'hf, 4'hc, 4'h0, 4'h3, 4'h3, 4'h1, 4'h4, 4'h5, 4'h3, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'hc, 4'h4, 4'h3, 4'hd, 4'hc, 4'h3, 4'h0, 4'h5, 4'h0, 4'h3, 4'h1, 4'hf, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0, 4'h5, 4'hc, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h4, 4'hc, 4'h4, 4'h0 };
assign dw_0[122] = dw_0_122[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_123 = { 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h7, 4'h3, 4'h3, 4'h1, 4'h1, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h7, 4'h4, 4'h3, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h3, 4'hc, 4'h0, 4'hf, 4'hc, 4'h5, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0 };
assign dw_0[123] = dw_0_123[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_124 = { 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h7, 4'h3, 4'h3, 4'h5, 4'h0, 4'hc, 4'hc, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h4, 4'h7, 4'hc, 4'hf, 4'h7, 4'h0, 4'hc, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'h0, 4'h3 };
assign dw_0[124] = dw_0_124[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_125 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h7, 4'h3, 4'hf, 4'h4, 4'h1, 4'hc, 4'hc, 4'h4, 4'h3, 4'h3, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'h5, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'h4, 4'h3 };
assign dw_0[125] = dw_0_125[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_126 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h7, 4'h3, 4'hf, 4'h4, 4'h3, 4'hc, 4'h3, 4'h0, 4'h3, 4'h7, 4'h4, 4'h4, 4'h5, 4'hc, 4'h0, 4'h3, 4'hf, 4'h0, 4'h4, 4'hc, 4'h5, 4'h4, 4'hc, 4'hc, 4'h4, 4'h3, 4'hd, 4'h0, 4'h3, 4'hc, 4'h4, 4'hc, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'h1, 4'h0, 4'hc, 4'h1, 4'hf, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h4, 4'hc, 4'h4, 4'h3 };
assign dw_0[126] = dw_0_126[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_127 = { 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'h7, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'hf, 4'h3, 4'h3, 4'h4, 4'h1, 4'h4, 4'h5, 4'h0, 4'h4, 4'hf, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'hf, 4'h7, 4'h0, 4'hd, 4'hd, 4'h0, 4'hc, 4'h5, 4'h0, 4'h1, 4'hc, 4'hf, 4'h5, 4'h0, 4'h1, 4'h0, 4'hc, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'hc, 4'h3, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0 };
assign dw_0[127] = dw_0_127[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_128 = { 4'h3, 4'h3, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h5, 4'h0, 4'hf, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'h1, 4'h1, 4'h0, 4'h5, 4'h3, 4'hf, 4'hd, 4'hc, 4'hd, 4'h0, 4'h4, 4'h4, 4'hf, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'hd, 4'h4, 4'hc, 4'hd, 4'hd, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h3, 4'hf, 4'hc, 4'hc, 4'hf, 4'h0, 4'h5, 4'h0, 4'h4, 4'hd, 4'h5, 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0 };
assign dw_0[128] = dw_0_128[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_129 = { 4'h1, 4'h1, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'h4, 4'hf, 4'h7, 4'hd, 4'h3, 4'hd, 4'h3, 4'hc, 4'h5, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'h1, 4'h0, 4'h7, 4'hc, 4'h3, 4'hd, 4'h4, 4'hc, 4'h0, 4'h4, 4'h4, 4'hf, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'hf, 4'h1, 4'h7, 4'h1, 4'h7, 4'h0, 4'h3, 4'h7, 4'h0, 4'h0 };
assign dw_0[129] = dw_0_129[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_130 = { 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'h7, 4'hf, 4'h3, 4'hc, 4'h3, 4'hd, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'h4, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'h1, 4'hf, 4'h5, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'hf, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h1, 4'hc, 4'h1, 4'h5, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0 };
assign dw_0[130] = dw_0_130[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_131 = { 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'hd, 4'h0, 4'hc, 4'h3, 4'hc, 4'h1, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h4, 4'hc, 4'hf, 4'hc, 4'hf, 4'h4, 4'h5, 4'hc, 4'h1, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h7, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[131] = dw_0_131[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_132 = { 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h4, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'hf, 4'hc, 4'h3, 4'h0, 4'h1, 4'h3, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4 };
assign dw_0[132] = dw_0_132[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_133 = { 4'h7, 4'hd, 4'hc, 4'h1, 4'h0, 4'hc, 4'h7, 4'h4, 4'hf, 4'h7, 4'hd, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'h7, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h7, 4'hf, 4'h3, 4'h5, 4'h0, 4'h3, 4'hd, 4'h7, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0 };
assign dw_0[133] = dw_0_133[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_134 = { 4'h4, 4'hc, 4'hc, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'hd, 4'hf, 4'hc, 4'hc, 4'h3, 4'h0, 4'h5, 4'h3, 4'h7, 4'hc, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h3, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'hf, 4'h5, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0 };
assign dw_0[134] = dw_0_134[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_135 = { 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h5, 4'h3, 4'h3, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'hc, 4'hc, 4'h4, 4'hc, 4'h0, 4'h3, 4'h1, 4'h1, 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'hf, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h1, 4'h3, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4 };
assign dw_0[135] = dw_0_135[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_136 = { 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'h4, 4'hf, 4'h0, 4'hd, 4'h0, 4'hd, 4'h7, 4'hd, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h7, 4'h0, 4'hf, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h7, 4'h3, 4'h3, 4'h5, 4'h1, 4'h1, 4'hc, 4'h7, 4'h4, 4'hf, 4'h3, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h4, 4'h4 };
assign dw_0[136] = dw_0_136[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_137 = { 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'hd, 4'hf, 4'h1, 4'hf, 4'hf, 4'h0, 4'h3, 4'h1, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h1, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3 };
assign dw_0[137] = dw_0_137[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_138 = { 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h5, 4'hc, 4'h3, 4'hc, 4'h3, 4'hc, 4'h3, 4'h0, 4'h4, 4'h7, 4'h1, 4'h0, 4'h3, 4'h7, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'hc, 4'h1, 4'h4, 4'h3, 4'hf, 4'h3, 4'h4, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'hf, 4'h3, 4'h0, 4'h4, 4'h0, 4'h7, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h1, 4'h4, 4'h0, 4'h7, 4'h0, 4'h7, 4'h0, 4'h4, 4'h3 };
assign dw_0[138] = dw_0_138[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_139 = { 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'hf, 4'h4, 4'h0, 4'h4, 4'h1, 4'h3, 4'hc, 4'h4, 4'h3, 4'h3, 4'h4, 4'h3, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'h7, 4'hc, 4'h3, 4'h1, 4'h0, 4'hd, 4'hc, 4'h4, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h5, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4 };
assign dw_0[139] = dw_0_139[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_140 = { 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h7, 4'h0, 4'h7, 4'hc, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'h5, 4'h4, 4'hc, 4'hd, 4'h7, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h1, 4'hf, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3 };
assign dw_0[140] = dw_0_140[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_141 = { 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h1, 4'h4, 4'hc, 4'h1, 4'h7, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'h3, 4'h3, 4'h1, 4'h0, 4'h1, 4'hc, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3 };
assign dw_0[141] = dw_0_141[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_142 = { 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'hc, 4'h4, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3, 4'hc, 4'h4, 4'h7, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'h7, 4'hc, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h7, 4'h4, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h7 };
assign dw_0[142] = dw_0_142[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_143 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h1, 4'h7, 4'h0, 4'h7, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'h3, 4'h5, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'hf, 4'h1, 4'hd, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h3, 4'h0, 4'h4, 4'h7, 4'h4, 4'h0 };
assign dw_0[143] = dw_0_143[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_144 = { 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h7, 4'h4, 4'hd, 4'hc, 4'h1, 4'h7, 4'h4, 4'h4, 4'h4, 4'h0, 4'h1, 4'hf, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h4, 4'h0, 4'hd, 4'h0, 4'h0, 4'h7, 4'hd, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h7, 4'h5, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h7, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0 };
assign dw_0[144] = dw_0_144[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_145 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h7, 4'h0, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'h7, 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h3, 4'h4, 4'hc, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h7, 4'h5, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'hc };
assign dw_0[145] = dw_0_145[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_146 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h3, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h7, 4'h3, 4'h1, 4'h0, 4'h3, 4'h1, 4'h0, 4'h5, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'h7, 4'h4, 4'h0, 4'h1, 4'h4, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h5, 4'hc, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[146] = dw_0_146[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_147 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h3, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h7, 4'h0, 4'h1, 4'h0, 4'h3, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h7, 4'h3, 4'h0, 4'h1, 4'h4, 4'h4, 4'h3, 4'h3, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h7, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h5, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[147] = dw_0_147[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_148 = { 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h7, 4'h0, 4'hd, 4'h3, 4'hd, 4'h0, 4'h4, 4'h4, 4'h7, 4'h0, 4'h1, 4'h7, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h7, 4'h7, 4'h3, 4'h1, 4'h0, 4'h4, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'h3, 4'h1, 4'hd, 4'h0, 4'h4, 4'hc, 4'hc, 4'h7, 4'h5, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[148] = dw_0_148[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_149 = { 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'hc, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'h7, 4'h0, 4'h1, 4'h7, 4'h3, 4'h3, 4'h4, 4'h1, 4'hc, 4'h0, 4'h1, 4'hc, 4'h0, 4'h4, 4'h1, 4'hd, 4'h0, 4'h0, 4'hc, 4'hc, 4'h4, 4'h5, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1 };
assign dw_0[149] = dw_0_149[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_150 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h4, 4'h1, 4'hd, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'h5, 4'hc, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1 };
assign dw_0[150] = dw_0_150[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_151 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'h1, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'h1, 4'h7, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h4, 4'h1, 4'hd, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0 };
assign dw_0[151] = dw_0_151[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_152 = { 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'hd, 4'h0, 4'hd, 4'h0, 4'h1, 4'h4, 4'h7, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'h7, 4'h3, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h1, 4'hc, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h5, 4'h3, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5 };
assign dw_0[152] = dw_0_152[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_153 = { 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h5, 4'h4, 4'h7, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'hc, 4'h1, 4'h7, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h4, 4'h5, 4'hf, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'h4 };
assign dw_0[153] = dw_0_153[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_154 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h3, 4'h3, 4'h1, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h7, 4'h0, 4'h1, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h7, 4'h0, 4'hd, 4'h4, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h4, 4'h5, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'hd, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0 };
assign dw_0[154] = dw_0_154[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_155 = { 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h7, 4'h3, 4'h1, 4'hd, 4'hd, 4'h0, 4'h0, 4'h4, 4'h7, 4'h0, 4'h1, 4'h3, 4'h3, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h7, 4'h7, 4'hf, 4'h1, 4'h4, 4'h7, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h5, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[155] = dw_0_155[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_156 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h7, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h7, 4'h0, 4'h1, 4'h4, 4'h3, 4'hd, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'hc, 4'h1, 4'h7, 4'h4, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'hc, 4'h0, 4'h4, 4'hf, 4'hc, 4'h4, 4'h4, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[156] = dw_0_156[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_157 = { 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h7, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h7, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'h3, 4'h1, 4'h4, 4'h1, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'hc, 4'h5, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0 };
assign dw_0[157] = dw_0_157[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_158 = { 4'h1, 4'h7, 4'hc, 4'h0, 4'h0, 4'h5, 4'h4, 4'h3, 4'h3, 4'hd, 4'hc, 4'h1, 4'h0, 4'h0, 4'h4, 4'h7, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'h3, 4'h4, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h4, 4'h5, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[158] = dw_0_158[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_159 = { 4'hd, 4'h3, 4'hc, 4'h0, 4'h0, 4'h5, 4'h5, 4'h7, 4'h3, 4'hd, 4'hf, 4'hd, 4'h4, 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'h5, 4'h0, 4'hd, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'h7, 4'h7, 4'h4, 4'h7, 4'hc, 4'h4, 4'hf, 4'h1, 4'h0, 4'h5, 4'h7, 4'h1, 4'hc, 4'h3, 4'hc, 4'hc, 4'hc, 4'h0, 4'h5, 4'h1, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'h4, 4'h5, 4'h0, 4'h1, 4'hf, 4'hc, 4'h0 };
assign dw_0[159] = dw_0_159[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_160 = { 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'h4, 4'h1, 4'h0, 4'h4, 4'h4, 4'hd, 4'h7, 4'h4, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h4, 4'hf, 4'h4, 4'hc, 4'h3, 4'hd, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h3, 4'h4, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc };
assign dw_0[160] = dw_0_160[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_161 = { 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h5, 4'hc, 4'h3, 4'h5, 4'h0, 4'hc, 4'hf, 4'h7, 4'h0, 4'hd, 4'hc, 4'h4, 4'h4, 4'hc, 4'hc, 4'h0, 4'h7, 4'hc, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf };
assign dw_0[161] = dw_0_161[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_162 = { 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'hd, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hc, 4'h3, 4'hd, 4'h0, 4'h3, 4'hc, 4'h7, 4'h0, 4'hd, 4'hc, 4'h0, 4'h7, 4'hf, 4'h3, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hf };
assign dw_0[162] = dw_0_162[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_163 = { 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h1, 4'hc, 4'h5, 4'h4, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h4, 4'h4, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h5, 4'hc, 4'h3, 4'h1, 4'h0, 4'hf, 4'hc, 4'h7, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'hf, 4'h0, 4'h3, 4'h7, 4'hc, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf };
assign dw_0[163] = dw_0_163[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_164 = { 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'hd, 4'h3, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'hc, 4'hf, 4'h1, 4'h0, 4'hf, 4'hc, 4'h7, 4'h3, 4'hc, 4'h0, 4'h5, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'hc, 4'hf, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc };
assign dw_0[164] = dw_0_164[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_165 = { 4'h3, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h1, 4'h3, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'hf, 4'h5, 4'hf, 4'hf, 4'h1, 4'h0, 4'hf, 4'hf, 4'h7, 4'h0, 4'hd, 4'h0, 4'h1, 4'h4, 4'hc, 4'hf, 4'h0, 4'h4, 4'hc, 4'h3, 4'h3, 4'h0, 4'hd, 4'h0, 4'h3, 4'h4, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf };
assign dw_0[165] = dw_0_165[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_166 = { 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'h1, 4'h7, 4'hc, 4'h3, 4'h3, 4'h3, 4'h0, 4'hc, 4'h3, 4'hc, 4'h4, 4'h0, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'h1, 4'h3, 4'h5, 4'hf, 4'hf, 4'h1, 4'h0, 4'hf, 4'hf, 4'h3, 4'h3, 4'hd, 4'hc, 4'h5, 4'h4, 4'hf, 4'hc, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'hc };
assign dw_0[166] = dw_0_166[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_167 = { 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h1, 4'hc, 4'h0, 4'h4, 4'hd, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h1, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'hf, 4'hf, 4'h1, 4'h0, 4'hf, 4'hc, 4'h7, 4'h3, 4'hc, 4'h4, 4'h5, 4'h0, 4'hf, 4'h3, 4'h0, 4'h7, 4'hc, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf };
assign dw_0[167] = dw_0_167[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_168 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'hd, 4'h3, 4'hd, 4'h4, 4'hc, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h5, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h5, 4'hc, 4'h3, 4'h1, 4'h0, 4'h3, 4'hf, 4'h3, 4'h3, 4'hf, 4'h0, 4'h4, 4'h4, 4'hf, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h4, 4'hd, 4'h0, 4'h3, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc };
assign dw_0[168] = dw_0_168[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_169 = { 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h1, 4'h7, 4'hd, 4'h3, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h5, 4'hc, 4'hf, 4'h1, 4'h0, 4'hf, 4'hc, 4'h7, 4'h0, 4'hd, 4'h0, 4'h5, 4'h4, 4'hf, 4'hc, 4'h0, 4'h7, 4'hd, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h1, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc };
assign dw_0[169] = dw_0_169[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_170 = { 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'hc, 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h5, 4'h0, 4'hf, 4'h0, 4'h1, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hc, 4'hf, 4'h1, 4'h0, 4'hf, 4'hc, 4'h7, 4'h0, 4'hd, 4'h0, 4'h0, 4'h4, 4'hf, 4'hc, 4'h0, 4'h4, 4'hd, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'h1, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc };
assign dw_0[170] = dw_0_170[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_171 = { 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h3, 4'h5, 4'hc, 4'h3, 4'h1, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf };
assign dw_0[171] = dw_0_171[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_172 = { 4'h1, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h5, 4'hf, 4'h3, 4'h1, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'hd, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf };
assign dw_0[172] = dw_0_172[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_173 = { 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'hf, 4'h4, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h4, 4'h1, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'hf, 4'h1, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'hc, 4'h0, 4'h1, 4'h4, 4'hc, 4'hc, 4'h0, 4'h4, 4'hc, 4'h3, 4'h3, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc };
assign dw_0[173] = dw_0_173[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_174 = { 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'h5, 4'hf, 4'h3, 4'h1, 4'h3, 4'hf, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'hf, 4'hc, 4'h0, 4'h3, 4'hd, 4'h0, 4'hc, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf };
assign dw_0[174] = dw_0_174[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_175 = { 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'hf, 4'h3, 4'h1, 4'h0, 4'h1, 4'h4, 4'hd, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'h3, 4'h1, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'hf, 4'h0, 4'h3, 4'h3, 4'hd, 4'h0, 4'hf, 4'h7, 4'hd, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc };
assign dw_0[175] = dw_0_175[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_176 = { 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h1, 4'hd, 4'h1, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'hd, 4'hf, 4'h3, 4'hc, 4'h0, 4'h3, 4'h7, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'h7, 4'h3, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h7, 4'h4, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[176] = dw_0_176[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_177 = { 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h1, 4'h1, 4'hd, 4'h1, 4'h3, 4'h0, 4'hd, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hc, 4'h0, 4'hf, 4'hd, 4'hc, 4'h7, 4'h0, 4'h4, 4'h0, 4'hf, 4'h4, 4'h3, 4'h1, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h3, 4'hd, 4'h0, 4'hd, 4'h0, 4'h0, 4'h7, 4'h4, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[177] = dw_0_177[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_178 = { 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'hd, 4'h1, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'hc, 4'h3, 4'hd, 4'h0, 4'hf, 4'h1, 4'h5, 4'h0, 4'hf, 4'h0, 4'h3, 4'h5, 4'h4, 4'hf, 4'h0, 4'h7, 4'h0, 4'h3, 4'hd, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h7, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0 };
assign dw_0[178] = dw_0_178[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_179 = { 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'hc, 4'hc, 4'hc, 4'h1, 4'h3, 4'h0, 4'h0, 4'h3, 4'h7, 4'h0, 4'h1, 4'hd, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hd, 4'hc, 4'h0, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'hf, 4'h4, 4'hf, 4'h1, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h3, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'hc, 4'h4 };
assign dw_0[179] = dw_0_179[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_180 = { 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'h3, 4'h4, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'hc, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h0, 4'hd, 4'h4, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[180] = dw_0_180[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_181 = { 4'h3, 4'hd, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'hc, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'hf, 4'h0, 4'h7, 4'h0, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[181] = dw_0_181[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_182 = { 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'hc, 4'hf, 4'hd, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h3, 4'h1, 4'h3, 4'h1, 4'h0, 4'h0, 4'h7, 4'h7, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[182] = dw_0_182[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_183 = { 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hd, 4'h3, 4'h0, 4'h0, 4'hd, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h5, 4'hc, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0 };
assign dw_0[183] = dw_0_183[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_184 = { 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'hc, 4'h1, 4'h0, 4'hd, 4'h1, 4'h3, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h5, 4'h0, 4'hd, 4'h0, 4'h0, 4'h7, 4'h7, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[184] = dw_0_184[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_185 = { 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h1, 4'h3, 4'hd, 4'h1, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h7, 4'h3, 4'h3, 4'h5, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0 };
assign dw_0[185] = dw_0_185[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_186 = { 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hd, 4'h3, 4'hc, 4'h1, 4'h3, 4'hd, 4'h1, 4'h3, 4'h4, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'h3, 4'hf, 4'hd, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h3, 4'h1, 4'h0, 4'h1, 4'h7, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[186] = dw_0_186[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_187 = { 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'hd, 4'h0, 4'h3, 4'hc, 4'h1, 4'h3, 4'h0, 4'h1, 4'h3, 4'hd, 4'h1, 4'h3, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hd, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0 };
assign dw_0[187] = dw_0_187[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_188 = { 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'hc, 4'hf, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hd, 4'h1, 4'h3, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'hd, 4'h3, 4'h3, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'hc, 4'hf, 4'h0, 4'h7, 4'h0, 4'h0, 4'h5, 4'h0, 4'hd, 4'h0, 4'h0, 4'h7, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[188] = dw_0_188[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_189 = { 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'h4, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h3, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[189] = dw_0_189[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_190 = { 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'hf, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'hd, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h3, 4'h1, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0 };
assign dw_0[190] = dw_0_190[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_191 = { 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1, 4'hd, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'h5, 4'hc, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0 };
assign dw_0[191] = dw_0_191[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_192 = { 4'h1, 4'hf, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h5, 4'h0, 4'h5, 4'h3, 4'h7, 4'h3, 4'h0, 4'hc, 4'h1, 4'h1, 4'h3, 4'h1, 4'h4, 4'h3, 4'hf, 4'h0, 4'h3, 4'h3, 4'h4, 4'h4, 4'h5, 4'h1, 4'h0, 4'hd, 4'h0, 4'hc, 4'hf, 4'h4, 4'h7, 4'h3, 4'h4, 4'h7, 4'hc, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'h4, 4'h1, 4'h3, 4'h4, 4'hf, 4'h1, 4'h0, 4'h7, 4'h4, 4'h0, 4'hd };
assign dw_0[192] = dw_0_192[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_193 = { 4'h1, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'hd, 4'h4, 4'h0, 4'h3, 4'h4, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h4, 4'h4, 4'h3, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h5, 4'h3, 4'h1, 4'h0, 4'hf, 4'h3, 4'hd, 4'h4, 4'h3, 4'h5, 4'h4, 4'h0, 4'hc, 4'h1, 4'h4, 4'h4, 4'h3, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd };
assign dw_0[193] = dw_0_193[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_194 = { 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'hf, 4'h4, 4'h4, 4'h3, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h1, 4'h3, 4'hd, 4'h0, 4'hf, 4'h0, 4'hc, 4'h4, 4'hf, 4'h4, 4'h4, 4'hc, 4'hc, 4'h1, 4'h7, 4'h4, 4'h3, 4'h3, 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'hf, 4'h1, 4'h0, 4'h4, 4'h0, 4'h4, 4'hc };
assign dw_0[194] = dw_0_194[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_195 = { 4'h1, 4'h5, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'hc, 4'h1, 4'h3, 4'h3, 4'hf, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'hd, 4'h0, 4'hf, 4'h1, 4'hc, 4'h4, 4'h3, 4'h4, 4'h3, 4'h0, 4'h3, 4'h1, 4'h4, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h7, 4'h3, 4'hd, 4'h0, 4'h1, 4'h0, 4'h3, 4'h1, 4'hc, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'hc };
assign dw_0[195] = dw_0_195[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_196 = { 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'h4, 4'h1, 4'h0, 4'hc, 4'h3, 4'h4, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'h3, 4'h4, 4'hf, 4'h3, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'hf, 4'h1, 4'hc, 4'h4, 4'h3, 4'h1, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'hc };
assign dw_0[196] = dw_0_196[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_197 = { 4'h1, 4'hc, 4'h4, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'h4, 4'h7, 4'h0, 4'h4, 4'h3, 4'h3, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'h7, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc };
assign dw_0[197] = dw_0_197[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_198 = { 4'hd, 4'hc, 4'h4, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'hd, 4'h0, 4'hd, 4'h3, 4'h0, 4'hf, 4'hf, 4'hc, 4'h1, 4'h0, 4'hc, 4'hf, 4'h4, 4'h3, 4'h3, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'hd, 4'h0, 4'hd, 4'h1, 4'hc, 4'h4, 4'h3, 4'h1, 4'hc, 4'hc, 4'h3, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h1, 4'h3, 4'h0, 4'h7, 4'hf, 4'h4, 4'hf };
assign dw_0[198] = dw_0_198[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_199 = { 4'h1, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'h1, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h5, 4'h4, 4'h3, 4'hd, 4'h3, 4'h0, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'hc };
assign dw_0[199] = dw_0_199[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_200 = { 4'hd, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'h1, 4'h1, 4'h0, 4'h4, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'hc, 4'h1, 4'hf, 4'h4, 4'hf, 4'h1, 4'h0, 4'hc, 4'hc, 4'hd, 4'h4, 4'h4, 4'h0, 4'h0, 4'h3, 4'hc, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'hc, 4'h0, 4'hc };
assign dw_0[200] = dw_0_200[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_201 = { 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h1, 4'h0, 4'hc, 4'hc, 4'h4, 4'h7, 4'hf, 4'h4, 4'hf, 4'h3, 4'h4, 4'h0, 4'h5, 4'hd, 4'hc, 4'h1, 4'h0, 4'hf, 4'h1, 4'hc, 4'h4, 4'h3, 4'h5, 4'h0, 4'h0, 4'hc, 4'hd, 4'h4, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'hc };
assign dw_0[201] = dw_0_201[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_202 = { 4'h1, 4'h0, 4'h4, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'h0, 4'h7, 4'h3, 4'h4, 4'h0, 4'hf, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h3, 4'h1, 4'hc, 4'h4, 4'h3, 4'h5, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'h5, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'hf };
assign dw_0[202] = dw_0_202[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_203 = { 4'hd, 4'h0, 4'h4, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'hf, 4'hf, 4'hc, 4'h1, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'hf, 4'hc, 4'h3, 4'h3, 4'h4, 4'h0, 4'h1, 4'h1, 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h7, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3, 4'hd, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'hc, 4'h1, 4'h0, 4'h4, 4'hc, 4'h0, 4'hc };
assign dw_0[203] = dw_0_203[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_204 = { 4'h1, 4'h1, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'hd, 4'h0, 4'hc, 4'h4, 4'h3, 4'h0, 4'h7, 4'hc, 4'hc, 4'h1, 4'h4, 4'h4, 4'h3, 4'h7, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'h4, 4'hc };
assign dw_0[204] = dw_0_204[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_205 = { 4'h1, 4'hd, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'h5, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h3, 4'h3, 4'h3, 4'h5, 4'h0, 4'hc, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'hd, 4'hc, 4'hc, 4'h3, 4'hd, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h4, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h4, 4'hd };
assign dw_0[205] = dw_0_205[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_206 = { 4'hd, 4'hd, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'h3, 4'h4, 4'h3, 4'h4, 4'hf, 4'hc, 4'h0, 4'h1, 4'h3, 4'h3, 4'h3, 4'h4, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h1, 4'h5, 4'h4, 4'h1, 4'hc, 4'hf, 4'h3, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h4, 4'hc, 4'h0, 4'h0, 4'h7, 4'h0, 4'h4, 4'hc };
assign dw_0[206] = dw_0_206[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_207 = { 4'h1, 4'hc, 4'h4, 4'h3, 4'h0, 4'hc, 4'hf, 4'h1, 4'hd, 4'h0, 4'h5, 4'h0, 4'h4, 4'hf, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h3, 4'h4, 4'h7, 4'h3, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'hf, 4'h3, 4'hc, 4'h4, 4'h3, 4'h4, 4'h5, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h3, 4'h7, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h4, 4'hc, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'hd };
assign dw_0[207] = dw_0_207[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_208 = { 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h7, 4'h4, 4'hf, 4'hc, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'h7, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'hd, 4'hc, 4'h0, 4'h7, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h3, 4'h7, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h4 };
assign dw_0[208] = dw_0_208[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_209 = { 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'h3, 4'h0, 4'h3, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'hd, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3 };
assign dw_0[209] = dw_0_209[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_210 = { 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'hf, 4'h0, 4'h3, 4'h4, 4'h3, 4'hc, 4'hc, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h7, 4'h5, 4'h7, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'hc, 4'h3, 4'h0, 4'hd, 4'h0, 4'h1, 4'hc, 4'h3, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h3 };
assign dw_0[210] = dw_0_210[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_211 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'hc, 4'h3, 4'h4, 4'h0, 4'hc, 4'hf, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h4, 4'hc, 4'h3, 4'h5, 4'h4, 4'h0, 4'h1, 4'h1, 4'hc, 4'h3, 4'hd, 4'h0, 4'hc, 4'h0, 4'h3, 4'h1, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h3, 4'h4, 4'h4 };
assign dw_0[211] = dw_0_211[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_212 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc, 4'hd, 4'h0, 4'hc, 4'h0, 4'h3, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'hc, 4'hf, 4'h7, 4'h0, 4'h0, 4'hd, 4'hc, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'h4, 4'h3 };
assign dw_0[212] = dw_0_212[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_213 = { 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'hf, 4'h0, 4'h3, 4'h4, 4'hf, 4'hc, 4'hc, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h4, 4'hd, 4'h7, 4'h0, 4'h7, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'hf, 4'h0, 4'h3, 4'hd, 4'h0, 4'h1, 4'h3, 4'h3, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h3 };
assign dw_0[213] = dw_0_213[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_214 = { 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'h4, 4'h3, 4'hd, 4'hc, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h7, 4'h5, 4'h7, 4'h0, 4'h0, 4'h0, 4'hd, 4'hf, 4'h1, 4'h0, 4'hc, 4'h4, 4'h7, 4'hd, 4'h0, 4'h1, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3 };
assign dw_0[214] = dw_0_214[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_215 = { 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h3, 4'h3, 4'h3, 4'h3, 4'h4, 4'h7, 4'hc, 4'hf, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'hd, 4'h7, 4'h4, 4'h3, 4'h0, 4'h1, 4'h0, 4'hd, 4'hc, 4'h1, 4'hc, 4'hc, 4'h0, 4'h4, 4'h1, 4'h0, 4'hd, 4'h0, 4'hf, 4'hc, 4'hc, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0 };
assign dw_0[215] = dw_0_215[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_216 = { 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h3, 4'hc, 4'hc, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'h4, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h4, 4'h4, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h4, 4'h3 };
assign dw_0[216] = dw_0_216[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_217 = { 4'h0, 4'h7, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h4, 4'h3, 4'hc, 4'hf, 4'h0, 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h1, 4'hf, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3 };
assign dw_0[217] = dw_0_217[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_218 = { 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h7, 4'h4, 4'h4, 4'h0, 4'h3, 4'h3, 4'hc, 4'h4, 4'h0, 4'hc, 4'hf, 4'h0, 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h4, 4'hc, 4'h3, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc, 4'h1, 4'hc, 4'hf, 4'h3, 4'h0, 4'h1, 4'h0, 4'hd, 4'h3, 4'h3, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3 };
assign dw_0[218] = dw_0_218[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_219 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'hf, 4'h0, 4'hc, 4'h4, 4'h0, 4'hd, 4'h3, 4'h0, 4'h3, 4'h7, 4'h0, 4'h0, 4'h4, 4'hf, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'hc, 4'h4, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0 };
assign dw_0[219] = dw_0_219[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_220 = { 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h4, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'hc, 4'h7, 4'h0, 4'h7, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h3, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0 };
assign dw_0[220] = dw_0_220[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_221 = { 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'hc, 4'h3, 4'h3, 4'hd, 4'h0, 4'hd, 4'h3, 4'h0, 4'h3, 4'hc, 4'h7, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3 };
assign dw_0[221] = dw_0_221[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_222 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'h4, 4'h3, 4'hc, 4'hc, 4'h0, 4'h3, 4'h7, 4'h3, 4'h4, 4'h4, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'hf, 4'h0, 4'h1, 4'h7, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0, 4'h3, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h7 };
assign dw_0[222] = dw_0_222[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_223 = { 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'h3, 4'h3, 4'hf, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h5, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'hc, 4'hd, 4'hd, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h3, 4'hc, 4'hf, 4'h7, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h3, 4'h4, 4'h7 };
assign dw_0[223] = dw_0_223[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_224 = { 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h1, 4'h3, 4'h0, 4'hd, 4'h1, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'hd, 4'h1, 4'hc, 4'hc, 4'h4, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h7, 4'h4, 4'h7, 4'h0, 4'hc, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h7, 4'h1, 4'h1, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3 };
assign dw_0[224] = dw_0_224[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_225 = { 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'hc, 4'hd, 4'h0, 4'h3, 4'hd, 4'h4, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc, 4'h4, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h1, 4'h0, 4'h4, 4'h4, 4'h4, 4'hc, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'hf };
assign dw_0[225] = dw_0_225[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_226 = { 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hd, 4'h1, 4'hf, 4'h0, 4'h1, 4'h1, 4'h7, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h4, 4'h7, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'h0 };
assign dw_0[226] = dw_0_226[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_227 = { 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h1, 4'hf, 4'hf, 4'h1, 4'hf, 4'h4, 4'h1, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'hc, 4'hd, 4'hc, 4'h4, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h5, 4'h3, 4'hc, 4'h0, 4'h4, 4'h3, 4'h3, 4'hc, 4'h4, 4'h4, 4'h4, 4'h0, 4'h4, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'hc };
assign dw_0[227] = dw_0_227[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_228 = { 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h4, 4'h0, 4'h7, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h7, 4'hc, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h3, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0 };
assign dw_0[228] = dw_0_228[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_229 = { 4'hd, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'hd, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h4, 4'h0, 4'h7, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0 };
assign dw_0[229] = dw_0_229[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_230 = { 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h3, 4'h0, 4'h4, 4'h1, 4'h7, 4'h1, 4'h7, 4'hf, 4'h3, 4'h3, 4'h3, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h4, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h3, 4'h1, 4'h0, 4'hd, 4'h0, 4'h4, 4'h1 };
assign dw_0[230] = dw_0_230[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_231 = { 4'hd, 4'hc, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'hc, 4'h5, 4'hc, 4'h7, 4'hd, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h7, 4'h0, 4'h4, 4'h0, 4'h5, 4'h7, 4'h1, 4'h3, 4'h0, 4'hc, 4'h3, 4'hc, 4'h4, 4'h4, 4'h4, 4'h4, 4'h4, 4'hc, 4'h1, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'hd };
assign dw_0[231] = dw_0_231[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_232 = { 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h4, 4'hc, 4'h4, 4'hd, 4'h4, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'hc, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h7, 4'hc, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'hf, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h1 };
assign dw_0[232] = dw_0_232[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_233 = { 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h7, 4'h1, 4'h4, 4'h3, 4'hf, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h3, 4'hd, 4'h0, 4'h1, 4'h3, 4'h3, 4'hc, 4'h4, 4'h4, 4'h7, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h7, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h1 };
assign dw_0[233] = dw_0_233[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_234 = { 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'h7, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'h4, 4'h3, 4'h3, 4'h1, 4'h0, 4'hc, 4'hd, 4'hc, 4'hc, 4'h0, 4'h4, 4'hc, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'hf, 4'h3, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0 };
assign dw_0[234] = dw_0_234[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_235 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h7, 4'hc, 4'h0, 4'hc, 4'h3, 4'h1, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h4, 4'h7, 4'hc, 4'h3, 4'h1, 4'hf, 4'h3, 4'h4, 4'h4, 4'h3, 4'h4, 4'hc, 4'h4, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0 };
assign dw_0[235] = dw_0_235[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_236 = { 4'hd, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hd, 4'h1, 4'hf, 4'hc, 4'h1, 4'h0, 4'h4, 4'h1, 4'h4, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h4, 4'h7, 4'hc, 4'h3, 4'h5, 4'hc, 4'h3, 4'hc, 4'h4, 4'h4, 4'h7, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h5, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h4, 4'h0 };
assign dw_0[236] = dw_0_236[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_237 = { 4'hd, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'hf, 4'hc, 4'h1, 4'hc, 4'h7, 4'hc, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h7, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h5, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0 };
assign dw_0[237] = dw_0_237[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_238 = { 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'h1, 4'hf, 4'hc, 4'h1, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h4, 4'h0, 4'h4, 4'h4, 4'hc, 4'h1, 4'h4, 4'hc, 4'h1, 4'hd, 4'h4, 4'h4, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'hf };
assign dw_0[238] = dw_0_238[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_239 = { 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'hf, 4'hc, 4'hd, 4'h3, 4'h0, 4'hd, 4'h4, 4'h0, 4'h3, 4'h3, 4'hd, 4'hf, 4'hd, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h4, 4'hc, 4'h4, 4'h4, 4'h1, 4'h0, 4'h1, 4'hc, 4'h1, 4'hc, 4'h3, 4'h7, 4'h1, 4'hd, 4'h4, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h1, 4'h1, 4'h7, 4'h0, 4'hd, 4'h0, 4'h0, 4'hf };
assign dw_0[239] = dw_0_239[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_240 = { 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h5, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h4, 4'h7, 4'hd, 4'h4, 4'hc, 4'h0, 4'hf, 4'h4, 4'h0, 4'hc, 4'h4, 4'h4, 4'h1, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0 };
assign dw_0[240] = dw_0_240[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_241 = { 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h7, 4'h1, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'hd, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'hf, 4'h0, 4'h0, 4'h4, 4'h3, 4'h1, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3, 4'hd, 4'h4, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'hc, 4'h0 };
assign dw_0[241] = dw_0_241[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_242 = { 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'h3, 4'h7, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h3, 4'h4, 4'h7, 4'h0, 4'hd, 4'h0, 4'h0, 4'h5, 4'h3, 4'h4, 4'h0, 4'h4, 4'h5, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[242] = dw_0_242[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_243 = { 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hd, 4'h1, 4'hc, 4'h1, 4'h3, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[243] = dw_0_243[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_244 = { 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'hf, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'hd, 4'h1, 4'h0, 4'h1, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h7, 4'h0, 4'h0, 4'h5, 4'h7, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0 };
assign dw_0[244] = dw_0_244[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_245 = { 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'hd, 4'h1, 4'hc, 4'h0, 4'h3, 4'h4, 4'hf, 4'h3, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0 };
assign dw_0[245] = dw_0_245[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_246 = { 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'hc, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'h4, 4'h1, 4'h1, 4'h4, 4'h4, 4'h1, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[246] = dw_0_246[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_247 = { 4'h4, 4'h3, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'hd, 4'h1, 4'hc, 4'h0, 4'hc, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'hf, 4'h4, 4'h1, 4'h0, 4'h4, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0 };
assign dw_0[247] = dw_0_247[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_248 = { 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'hf, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[248] = dw_0_248[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_249 = { 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h7, 4'h0, 4'hf, 4'h3, 4'h4, 4'h1, 4'hf, 4'hc, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'h0, 4'h1, 4'h4, 4'hd, 4'h1, 4'h3, 4'h4, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0 };
assign dw_0[249] = dw_0_249[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_250 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'hd, 4'h0, 4'hc, 4'h7, 4'h0, 4'hd, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0 };
assign dw_0[250] = dw_0_250[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_251 = { 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h5, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h4, 4'h7, 4'h3, 4'h0, 4'h4, 4'hc, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'hf, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[251] = dw_0_251[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_252 = { 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hd, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0 };
assign dw_0[252] = dw_0_252[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_253 = { 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h3, 4'h4, 4'hc, 4'h0, 4'h7, 4'h1, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'hd, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3 };
assign dw_0[253] = dw_0_253[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_254 = { 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h5, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[254] = dw_0_254[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_255 = { 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'h0, 4'h4, 4'hd, 4'h3, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h7, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h4, 4'h4, 4'hc, 4'hf, 4'hc, 4'h0, 4'h1, 4'hf, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[255] = dw_0_255[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_256 = { 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'h3, 4'h0, 4'h4, 4'h4, 4'h7, 4'h0, 4'h1, 4'h1, 4'hc, 4'hc, 4'hc, 4'h4, 4'h1, 4'h7, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h1, 4'h1, 4'h3, 4'h0, 4'h1, 4'hf, 4'h0, 4'hd, 4'h4, 4'hd, 4'h0, 4'h4, 4'h4, 4'hc, 4'h0 };
assign dw_0[256] = dw_0_256[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_257 = { 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'h7, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'hf, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'h4, 4'h0, 4'h3, 4'h7, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h7, 4'h1, 4'h0, 4'h4, 4'h4, 4'hc, 4'h4 };
assign dw_0[257] = dw_0_257[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_258 = { 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h4, 4'hc, 4'h0, 4'h3, 4'hc, 4'h4, 4'h4, 4'h1, 4'h4, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'h1, 4'h0, 4'hf, 4'h0, 4'h1, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hd, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1 };
assign dw_0[258] = dw_0_258[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_259 = { 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h5, 4'h4, 4'h1, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h4, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'h1, 4'h3, 4'h4, 4'h1, 4'h3, 4'h0, 4'hd, 4'h5, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5 };
assign dw_0[259] = dw_0_259[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_260 = { 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h1, 4'h3, 4'h0, 4'h5, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h4, 4'h1, 4'h3, 4'h0, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1 };
assign dw_0[260] = dw_0_260[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_261 = { 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'hc, 4'h3, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h7, 4'h5, 4'hc, 4'h1, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hd, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'hd, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1 };
assign dw_0[261] = dw_0_261[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_262 = { 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'hc, 4'h3, 4'h5, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h7, 4'h1, 4'h0, 4'h1, 4'h3, 4'h3, 4'h5, 4'h7, 4'hd, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[262] = dw_0_262[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_263 = { 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h7, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h7, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h1, 4'hf, 4'h4, 4'h0, 4'h3, 4'h4, 4'h1, 4'h5, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1 };
assign dw_0[263] = dw_0_263[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_264 = { 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h7, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'hc, 4'h4, 4'hd, 4'h7, 4'hc, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h5, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h7, 4'hc, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1 };
assign dw_0[264] = dw_0_264[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_265 = { 4'h0, 4'h4, 4'hc, 4'h1, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h4, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h4, 4'h1, 4'h3, 4'h3, 4'h5, 4'h7, 4'hc, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5 };
assign dw_0[265] = dw_0_265[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_266 = { 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h4, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'hc, 4'h0, 4'hc, 4'h4, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h7, 4'hc, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'h7, 4'h3, 4'h0, 4'h1, 4'h1, 4'h3, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h5 };
assign dw_0[266] = dw_0_266[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_267 = { 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'hd, 4'h5, 4'h0, 4'h4, 4'h1, 4'hd, 4'h0, 4'hc, 4'h0, 4'h5, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h5, 4'h3, 4'h0, 4'h7, 4'h3, 4'h0, 4'h1, 4'h4, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1 };
assign dw_0[267] = dw_0_267[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_268 = { 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h1, 4'h0, 4'h3, 4'h3, 4'h5, 4'h3, 4'h0, 4'h7, 4'h3, 4'h4, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[268] = dw_0_268[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_269 = { 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'hd, 4'h4, 4'h1, 4'h7, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1 };
assign dw_0[269] = dw_0_269[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_270 = { 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'hd, 4'h4, 4'hc, 4'h4, 4'h0, 4'h1, 4'h3, 4'h3, 4'h0, 4'h1, 4'h3, 4'h1, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h7, 4'h5, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h1, 4'h7, 4'h1, 4'h0, 4'h7, 4'h0, 4'hc, 4'h5 };
assign dw_0[270] = dw_0_270[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_271 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h0, 4'h3, 4'hc, 4'h4, 4'h0, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'hc, 4'h0, 4'hc, 4'h4, 4'h1, 4'h3, 4'h0, 4'hd, 4'h3, 4'h3, 4'h0, 4'h1, 4'hf, 4'h0, 4'hc, 4'hc, 4'hc, 4'h1, 4'h0, 4'h1, 4'h4, 4'h7, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hf, 4'h7, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1 };
assign dw_0[271] = dw_0_271[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_272 = { 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'hc, 4'h4, 4'h7, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'hc, 4'hc, 4'h1, 4'hc, 4'h7, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hd, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'hc, 4'hc, 4'h1 };
assign dw_0[272] = dw_0_272[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_273 = { 4'hf, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'hd, 4'h0, 4'h3, 4'h4, 4'hf, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'hf, 4'hd, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hd, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0 };
assign dw_0[273] = dw_0_273[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_274 = { 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'h4, 4'h7, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h7, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h5, 4'hc, 4'hc, 4'hc, 4'hc, 4'h0, 4'h3, 4'h4, 4'hc, 4'h0, 4'hc, 4'h1, 4'hd, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0 };
assign dw_0[274] = dw_0_274[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_275 = { 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'hf, 4'hc, 4'h4, 4'h0, 4'h0, 4'hf, 4'h5, 4'hc, 4'hc, 4'hd, 4'hc, 4'h4, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[275] = dw_0_275[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_276 = { 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h4, 4'h4, 4'h4, 4'h4, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'hc, 4'hd, 4'hc, 4'h4, 4'h3, 4'h4, 4'hc, 4'h0, 4'h1, 4'h3, 4'hd, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'hd, 4'h0, 4'h0 };
assign dw_0[276] = dw_0_276[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_277 = { 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'h1, 4'hf, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h4, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hd, 4'h5, 4'hc, 4'hc, 4'h1, 4'hc, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0 };
assign dw_0[277] = dw_0_277[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_278 = { 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'hc, 4'hc, 4'h4, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h1, 4'h3, 4'h3, 4'h3, 4'h5, 4'hc, 4'hc, 4'h1, 4'hc, 4'h1, 4'h1, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h1 };
assign dw_0[278] = dw_0_278[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_279 = { 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hc, 4'h5, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h4, 4'hc, 4'h0, 4'hc, 4'hc, 4'hd, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0 };
assign dw_0[279] = dw_0_279[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_280 = { 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'hd, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h5, 4'hc, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h7, 4'h0, 4'h0, 4'h3, 4'hc, 4'hd, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h1 };
assign dw_0[280] = dw_0_280[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_281 = { 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'hf, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h5, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0 };
assign dw_0[281] = dw_0_281[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_282 = { 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h5, 4'h3, 4'h0, 4'h4, 4'h1, 4'hc, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h7, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'hc, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'hc, 4'h0, 4'hd, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[282] = dw_0_282[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_283 = { 4'h3, 4'h7, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h7, 4'h1, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0, 4'hd, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0 };
assign dw_0[283] = dw_0_283[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_284 = { 4'hf, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h7, 4'h1, 4'hc, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h5, 4'h3, 4'h0, 4'h0, 4'h5, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h4, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'hd, 4'hc, 4'hc, 4'hc };
assign dw_0[284] = dw_0_284[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_285 = { 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'h4, 4'hd, 4'hc, 4'h0, 4'h1, 4'h3, 4'hc, 4'h1, 4'h3, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'hf, 4'hd, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h5, 4'h0, 4'hc, 4'h4, 4'hf, 4'hd, 4'h3, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0 };
assign dw_0[285] = dw_0_285[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_286 = { 4'hf, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'hd, 4'h0, 4'h4, 4'h5, 4'h0, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'hd, 4'hc, 4'h0, 4'hc };
assign dw_0[286] = dw_0_286[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_287 = { 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h3, 4'hd, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0 };
assign dw_0[287] = dw_0_287[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_288 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'hf, 4'hc, 4'h3, 4'h1, 4'hc, 4'h5, 4'h4, 4'h0, 4'h3, 4'h3, 4'h7, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'h5, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'hf, 4'h0, 4'h0, 4'hd, 4'h3, 4'hd, 4'hd, 4'h4, 4'h4, 4'h0, 4'h7, 4'hd, 4'h1, 4'h1, 4'h1, 4'h4, 4'h0, 4'h1, 4'h5, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0 };
assign dw_0[288] = dw_0_288[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_289 = { 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h4, 4'h7, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'hc, 4'h5, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h5, 4'hc, 4'h4, 4'h4, 4'h4, 4'h3, 4'hd, 4'hf, 4'h7, 4'h3, 4'h4, 4'hf, 4'h1, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h3, 4'h4, 4'hc, 4'h0, 4'h0, 4'hd, 4'h4, 4'h1 };
assign dw_0[289] = dw_0_289[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_290 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'hc, 4'h5, 4'h7, 4'h0, 4'h0, 4'h1, 4'h4, 4'h3, 4'h3, 4'h0, 4'h4, 4'hc, 4'h1, 4'h5, 4'hc, 4'h0, 4'h7, 4'h4, 4'h0, 4'hd, 4'h3, 4'h4, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc, 4'h4, 4'h4, 4'h0, 4'h3, 4'hd, 4'h5, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0, 4'h1, 4'h1, 4'hf, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'h4 };
assign dw_0[290] = dw_0_290[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_291 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h1, 4'h3, 4'h5, 4'hc, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1, 4'h5, 4'hc, 4'h0, 4'h4, 4'h4, 4'h3, 4'h1, 4'hf, 4'h3, 4'h0, 4'h4, 4'h0, 4'h1, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h1, 4'h1, 4'h4, 4'h3, 4'h1, 4'h7, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h5, 4'h4, 4'h5 };
assign dw_0[291] = dw_0_291[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_292 = { 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'hc, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h7, 4'h3, 4'h1, 4'h3, 4'h1, 4'hc, 4'h1, 4'h5, 4'h0, 4'h0, 4'h3, 4'h7, 4'h0, 4'h0, 4'hf, 4'h7, 4'h0, 4'h4, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h5, 4'h0, 4'hd, 4'h0, 4'h4, 4'h3, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5 };
assign dw_0[292] = dw_0_292[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_293 = { 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h1, 4'hc, 4'h5, 4'h4, 4'h0, 4'h3, 4'h1, 4'h7, 4'h1, 4'hc, 4'h0, 4'h5, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'hf, 4'h7, 4'h0, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h1, 4'h7, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h3, 4'h5, 4'h4, 4'h4 };
assign dw_0[293] = dw_0_293[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_294 = { 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'hf, 4'h1, 4'hc, 4'h5, 4'h3, 4'h1, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h5, 4'hc, 4'h0, 4'h4, 4'h4, 4'h3, 4'hc, 4'hf, 4'h7, 4'h1, 4'h5, 4'h3, 4'h1, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'hd, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h7, 4'h1, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'h3, 4'h4, 4'hc, 4'h0, 4'h3, 4'h1, 4'h4, 4'h5 };
assign dw_0[294] = dw_0_294[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_295 = { 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'h5, 4'hc, 4'h0, 4'h4, 4'h4, 4'h3, 4'hc, 4'hf, 4'h7, 4'h0, 4'h5, 4'h0, 4'hd, 4'h1, 4'h0, 4'h0, 4'h1, 4'h7, 4'hd, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'hd, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1 };
assign dw_0[295] = dw_0_295[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_296 = { 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'h5, 4'h0, 4'hd, 4'h3, 4'h1, 4'h7, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'h5, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'hf, 4'h4, 4'h1, 4'h3, 4'h3, 4'h1, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h4, 4'h4, 4'h1, 4'h7, 4'h4, 4'h0, 4'h0, 4'h5, 4'hf, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5 };
assign dw_0[296] = dw_0_296[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_297 = { 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h5, 4'h7, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'hc, 4'h0, 4'h7, 4'h7, 4'hf, 4'h0, 4'hf, 4'h7, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'hd, 4'h0, 4'h0, 4'h7, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'h5 };
assign dw_0[297] = dw_0_297[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_298 = { 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h5, 4'h7, 4'h3, 4'hc, 4'h0, 4'hf, 4'h1, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h7, 4'h0, 4'hd, 4'h3, 4'h4, 4'hc, 4'h1, 4'h5, 4'hc, 4'h0, 4'h7, 4'h4, 4'h3, 4'h0, 4'hf, 4'h7, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'h5 };
assign dw_0[298] = dw_0_298[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_299 = { 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h7, 4'h1, 4'h3, 4'hc, 4'h1, 4'h0, 4'h5, 4'h4, 4'h0, 4'hd, 4'h1, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h1, 4'h5, 4'hc, 4'h0, 4'h4, 4'h4, 4'hc, 4'h0, 4'hf, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5 };
assign dw_0[299] = dw_0_299[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_300 = { 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h7, 4'hd, 4'hc, 4'h0, 4'h1, 4'hc, 4'h5, 4'h0, 4'h1, 4'h0, 4'h1, 4'h7, 4'hc, 4'hc, 4'h0, 4'h4, 4'hc, 4'h1, 4'h5, 4'hc, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h5, 4'h7, 4'h0, 4'h3, 4'h1, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h5 };
assign dw_0[300] = dw_0_300[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_301 = { 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h1, 4'hc, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h7, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'h5, 4'hc, 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h5, 4'h7, 4'h0, 4'h3, 4'h1, 4'h5, 4'hc, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h1 };
assign dw_0[301] = dw_0_301[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_302 = { 4'h0, 4'h5, 4'hc, 4'h1, 4'h0, 4'h4, 4'h4, 4'h1, 4'hf, 4'h0, 4'h3, 4'h1, 4'hd, 4'h5, 4'h7, 4'h1, 4'h3, 4'h3, 4'h7, 4'h3, 4'h1, 4'hc, 4'h4, 4'hc, 4'h1, 4'h5, 4'hc, 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'hd, 4'h4, 4'h0, 4'h5, 4'h7, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h3, 4'h5, 4'h0, 4'h0, 4'hc, 4'h1, 4'h1, 4'hc, 4'h4, 4'h4, 4'h0, 4'h3, 4'hc, 4'h4, 4'h5 };
assign dw_0[302] = dw_0_302[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_303 = { 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h5, 4'h7, 4'h5, 4'hc, 4'hc, 4'h0, 4'h1, 4'hd, 4'h5, 4'h4, 4'hc, 4'h3, 4'h3, 4'h7, 4'h0, 4'h0, 4'hc, 4'h5, 4'hc, 4'h5, 4'h5, 4'hc, 4'h0, 4'h4, 4'h7, 4'h3, 4'h0, 4'hc, 4'h4, 4'h3, 4'h0, 4'h3, 4'hd, 4'hc, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h7, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h5 };
assign dw_0[303] = dw_0_303[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_304 = { 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'h5, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h1, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'hc, 4'hc, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0 };
assign dw_0[304] = dw_0_304[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_305 = { 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h1, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h1, 4'hf, 4'hc, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h3, 4'h5, 4'h0, 4'h0, 4'h5, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h3 };
assign dw_0[305] = dw_0_305[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_306 = { 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'hd, 4'h0, 4'h7, 4'h0, 4'h3, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3, 4'hc, 4'h1, 4'hc, 4'h0, 4'hc, 4'hd, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h4, 4'h7, 4'h4, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0 };
assign dw_0[306] = dw_0_306[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_307 = { 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h1, 4'h3, 4'h3, 4'h1, 4'hf, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h7, 4'h3, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'h1, 4'h3, 4'hc, 4'hf, 4'hd, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'hf, 4'hf, 4'h1, 4'h0, 4'h0, 4'h4, 4'h7, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[307] = dw_0_307[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_308 = { 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'hf, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hd, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h5, 4'h4, 4'h7, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3 };
assign dw_0[308] = dw_0_308[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_309 = { 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h1, 4'hf, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h3, 4'hf, 4'h3, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hd, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h1, 4'hf, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h5, 4'h7, 4'h7, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0 };
assign dw_0[309] = dw_0_309[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_310 = { 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h1, 4'h3, 4'h3, 4'h0, 4'h3, 4'h4, 4'hf, 4'hc, 4'hc, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'hf, 4'hc, 4'hf, 4'h3, 4'h3, 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0 };
assign dw_0[310] = dw_0_310[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_311 = { 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'h3, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'hc, 4'h1, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h0, 4'h3, 4'hf, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3 };
assign dw_0[311] = dw_0_311[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_312 = { 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h5, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'hf, 4'h3, 4'h3, 4'h1, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'hf, 4'hc, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'hc, 4'h1, 4'hf, 4'hc, 4'hf, 4'hc, 4'h3, 4'hc, 4'h0, 4'h7, 4'h3, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'h0, 4'h5, 4'h7, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'hc };
assign dw_0[312] = dw_0_312[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_313 = { 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hf, 4'h0, 4'hf, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h1, 4'h0, 4'hc, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc };
assign dw_0[313] = dw_0_313[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_314 = { 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'hc, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'hf, 4'hd, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'hc, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'h1, 4'h4, 4'h7, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf };
assign dw_0[314] = dw_0_314[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_315 = { 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'hf, 4'h1, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h4, 4'hd, 4'h0, 4'hd, 4'hc, 4'hc, 4'h1, 4'h3, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3 };
assign dw_0[315] = dw_0_315[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_316 = { 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h3, 4'h0, 4'h3, 4'h4, 4'hf, 4'hc, 4'hc, 4'h1, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'hc, 4'hc, 4'hc, 4'h1, 4'hc, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4, 4'hf, 4'h1, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h3 };
assign dw_0[316] = dw_0_316[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_317 = { 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hd, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h4, 4'h0, 4'h3, 4'h4, 4'h3, 4'h7, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h4, 4'h0, 4'hf, 4'hc, 4'h5, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h3, 4'h3, 4'h7, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0 };
assign dw_0[317] = dw_0_317[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_318 = { 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h7, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'hf, 4'h1, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h7, 4'h0, 4'h3, 4'hf, 4'h5, 4'h0, 4'h0, 4'h5, 4'h4, 4'h7, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3 };
assign dw_0[318] = dw_0_318[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_319 = { 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h7, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf };
assign dw_0[319] = dw_0_319[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_320 = { 4'h7, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'hf, 4'h5, 4'h4, 4'h3, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'hc, 4'hc, 4'hc, 4'hc, 4'h4, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h3, 4'h3, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0 };
assign dw_0[320] = dw_0_320[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_321 = { 4'h3, 4'h7, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'hc, 4'hc, 4'h7, 4'hf, 4'hc, 4'h7, 4'hd, 4'hc, 4'hf, 4'h1, 4'h1, 4'h1, 4'h5, 4'h3, 4'h4, 4'h3, 4'h4, 4'h7, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'h0, 4'h4, 4'h1, 4'h0, 4'h5, 4'hc, 4'hc, 4'hc, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'hd, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf };
assign dw_0[321] = dw_0_321[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_322 = { 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h1, 4'hf, 4'h7, 4'h3, 4'h3, 4'h4, 4'hd, 4'hc, 4'hc, 4'h0, 4'h0, 4'hd, 4'h1, 4'h3, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h7, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc };
assign dw_0[322] = dw_0_322[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_323 = { 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'h7, 4'h3, 4'h0, 4'h4, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'h7, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'hc, 4'h1, 4'hc, 4'hd, 4'h0, 4'hc, 4'h4, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'hf, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3 };
assign dw_0[323] = dw_0_323[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_324 = { 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h7, 4'h3, 4'h0, 4'h7, 4'h1, 4'hc, 4'hf, 4'h1, 4'h3, 4'hc, 4'h1, 4'h3, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hc, 4'h1, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h1, 4'h3, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'h4, 4'hc };
assign dw_0[324] = dw_0_324[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_325 = { 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h7, 4'h7, 4'h0, 4'h7, 4'hd, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h5, 4'h3, 4'h1, 4'h0, 4'h0, 4'h7, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h7, 4'h4, 4'h4, 4'h3, 4'h3, 4'hc, 4'h5, 4'hf, 4'hc, 4'h3, 4'hc, 4'h4, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h4, 4'hd, 4'h5, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'hf };
assign dw_0[325] = dw_0_325[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_326 = { 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h4, 4'h3, 4'hf, 4'h4, 4'hd, 4'hc, 4'hc, 4'h0, 4'h3, 4'h5, 4'h5, 4'h3, 4'h1, 4'h3, 4'h4, 4'h7, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hd, 4'h5, 4'hc, 4'hc, 4'h0, 4'hc, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'hd, 4'hd, 4'h3, 4'h4, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc };
assign dw_0[326] = dw_0_326[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_327 = { 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h7, 4'h3, 4'h3, 4'h4, 4'hd, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h3, 4'hc, 4'h5, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'hd, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0 };
assign dw_0[327] = dw_0_327[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_328 = { 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h4, 4'h3, 4'h3, 4'h4, 4'hd, 4'hc, 4'h3, 4'h1, 4'h3, 4'h1, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'hc, 4'h0, 4'hc, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h1, 4'hc, 4'hc, 4'h0, 4'hc, 4'h1, 4'hc, 4'h3, 4'h1, 4'h0, 4'h0, 4'h4, 4'hd, 4'hd, 4'h0, 4'h0, 4'h0, 4'h1, 4'hd, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc };
assign dw_0[328] = dw_0_328[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_329 = { 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h4, 4'hd, 4'hc, 4'h0, 4'h1, 4'h3, 4'hd, 4'h5, 4'h3, 4'h0, 4'h3, 4'h0, 4'h7, 4'hc, 4'hc, 4'h0, 4'hc, 4'hc, 4'h3, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'h5, 4'hc, 4'hc, 4'hc, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'hd, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0 };
assign dw_0[329] = dw_0_329[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_330 = { 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'h3, 4'h4, 4'h3, 4'h3, 4'h4, 4'h1, 4'hc, 4'h0, 4'h1, 4'h3, 4'h1, 4'h4, 4'h3, 4'h4, 4'h3, 4'h4, 4'h4, 4'h0, 4'hf, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'hd, 4'h1, 4'hc, 4'hd, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0 };
assign dw_0[330] = dw_0_330[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_331 = { 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hd, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'hd, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h5, 4'h3, 4'h4, 4'h3, 4'h4, 4'h7, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0 };
assign dw_0[331] = dw_0_331[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_332 = { 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'h3, 4'hf, 4'h4, 4'hd, 4'hc, 4'hf, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h7, 4'h3, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h4, 4'hf, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hd, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0 };
assign dw_0[332] = dw_0_332[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_333 = { 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h7, 4'h3, 4'h3, 4'h4, 4'hd, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'h7, 4'hf, 4'hc, 4'h0, 4'hf, 4'h0, 4'h7, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h1, 4'hc, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h3, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0 };
assign dw_0[333] = dw_0_333[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_334 = { 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'hc, 4'hf, 4'h4, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'h4, 4'h4, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h5, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc };
assign dw_0[334] = dw_0_334[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_335 = { 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'hd, 4'h4, 4'h3, 4'h3, 4'h4, 4'hd, 4'hc, 4'hc, 4'h1, 4'h1, 4'hd, 4'h1, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'hc, 4'h7, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h7, 4'hd, 4'h1, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc };
assign dw_0[335] = dw_0_335[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_336 = { 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h5, 4'h1, 4'hd, 4'h0, 4'h4, 4'h3, 4'h4, 4'h7, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h4, 4'h7, 4'h0, 4'h3, 4'hc, 4'h4, 4'h1, 4'h3, 4'h4, 4'hc, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'h1, 4'h4, 4'h4, 4'h7, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0 };
assign dw_0[336] = dw_0_336[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_337 = { 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'h3, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h7, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'hc, 4'hc, 4'h4, 4'hd, 4'h3, 4'h0, 4'hd, 4'h3, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h5, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc };
assign dw_0[337] = dw_0_337[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_338 = { 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'hd, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'h3, 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h3, 4'h3, 4'hd, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h7, 4'h1, 4'h0, 4'h4, 4'hc, 4'hc, 4'h0 };
assign dw_0[338] = dw_0_338[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_339 = { 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h7, 4'h3, 4'h0, 4'h1, 4'h7, 4'h1, 4'h3, 4'h3, 4'hd, 4'h0, 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'hd, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0 };
assign dw_0[339] = dw_0_339[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_340 = { 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h0, 4'h4, 4'hd, 4'h3, 4'h0, 4'hd, 4'h3, 4'hd, 4'h4, 4'hc, 4'h0, 4'h0, 4'hd, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h4, 4'h7, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0 };
assign dw_0[340] = dw_0_340[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_341 = { 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h7, 4'h3, 4'h3, 4'h3, 4'h3, 4'h1, 4'h0, 4'h1, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h7, 4'h4, 4'h0, 4'h4, 4'hd, 4'h3, 4'hc, 4'hd, 4'h3, 4'h0, 4'h5, 4'hc, 4'h5, 4'h4, 4'hd, 4'h4, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h7, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1 };
assign dw_0[341] = dw_0_341[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_342 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h1, 4'hd, 4'h1, 4'h0, 4'hd, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h3, 4'h3, 4'hd, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h5, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0 };
assign dw_0[342] = dw_0_342[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_343 = { 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4, 4'h1, 4'h3, 4'h3, 4'hd, 4'hf, 4'hd, 4'h4, 4'h0, 4'h4, 4'h1, 4'hd, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0 };
assign dw_0[343] = dw_0_343[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_344 = { 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'hc, 4'h4, 4'h3, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h7, 4'hd, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h5, 4'h0, 4'hc, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0 };
assign dw_0[344] = dw_0_344[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_345 = { 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'hc, 4'h7, 4'h0, 4'h1, 4'h3, 4'h1, 4'h0, 4'hc, 4'h4, 4'h7, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'h4, 4'hd, 4'h3, 4'h0, 4'hd, 4'hf, 4'h4, 4'h5, 4'h0, 4'h4, 4'h4, 4'hc, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1 };
assign dw_0[345] = dw_0_345[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_346 = { 4'h1, 4'h7, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'h3, 4'h1, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h1, 4'h7, 4'hd, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'h4, 4'h0, 4'hc, 4'hd, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[346] = dw_0_346[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_347 = { 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h5, 4'hd, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0 };
assign dw_0[347] = dw_0_347[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_348 = { 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'h0, 4'h4, 4'hd, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h3, 4'h3, 4'h3, 4'hc, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0 };
assign dw_0[348] = dw_0_348[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_349 = { 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h4, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0 };
assign dw_0[349] = dw_0_349[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_350 = { 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h7, 4'h7, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'hc, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0 };
assign dw_0[350] = dw_0_350[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_351 = { 4'h1, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h1, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'hd, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'h3, 4'h3, 4'hf, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h7, 4'h5, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0 };
assign dw_0[351] = dw_0_351[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_352 = { 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h4, 4'h0, 4'hd, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h1, 4'h0, 4'h7, 4'h0, 4'h7, 4'hc, 4'h4, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h4, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h4, 4'h0 };
assign dw_0[352] = dw_0_352[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_353 = { 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hd, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h1, 4'hf, 4'h7, 4'h0, 4'h4, 4'hc, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h7, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0 };
assign dw_0[353] = dw_0_353[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_354 = { 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h3, 4'h1, 4'hc, 4'h3, 4'h3, 4'h0, 4'hc, 4'h4, 4'h4, 4'h4, 4'hc, 4'h4, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[354] = dw_0_354[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_355 = { 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'h3, 4'h1, 4'h3, 4'h4, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h7, 4'h3, 4'h4, 4'hc, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h7, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'hc };
assign dw_0[355] = dw_0_355[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_356 = { 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h3, 4'hc, 4'h1, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h7, 4'h0, 4'h4, 4'hc, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'hc };
assign dw_0[356] = dw_0_356[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_357 = { 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h4, 4'h3, 4'hd, 4'h0, 4'hf, 4'h3, 4'h3, 4'hc, 4'h3, 4'h0, 4'h4, 4'hd, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h5, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'h0 };
assign dw_0[357] = dw_0_357[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_358 = { 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'h3, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h7, 4'h0, 4'h7, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h7, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0 };
assign dw_0[358] = dw_0_358[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_359 = { 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h5, 4'h3, 4'h4, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'h4, 4'h0, 4'h5, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h7, 4'h0, 4'h4, 4'hc, 4'h0, 4'hc, 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'h5, 4'h7, 4'h0, 4'hc, 4'hd, 4'h0, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0 };
assign dw_0[359] = dw_0_359[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_360 = { 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h1, 4'h3, 4'h1, 4'h3, 4'hc, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc, 4'h4, 4'hd, 4'h1, 4'hf, 4'h3, 4'h0, 4'h0, 4'h5, 4'h7, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h3, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0 };
assign dw_0[360] = dw_0_360[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_361 = { 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h3, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h3, 4'hf, 4'h3, 4'h3, 4'h0, 4'h7, 4'h4, 4'h4, 4'hd, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4, 4'h5, 4'h4, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'hf, 4'h4, 4'h3, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h1 };
assign dw_0[361] = dw_0_361[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_362 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h4, 4'hf, 4'h3, 4'h0, 4'hc, 4'h1, 4'hd, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'hc, 4'hc, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0 };
assign dw_0[362] = dw_0_362[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_363 = { 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'hc, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h1, 4'h4, 4'hd, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'h5, 4'h7, 4'h0, 4'hc, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0 };
assign dw_0[363] = dw_0_363[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_364 = { 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h7, 4'h3, 4'h1, 4'h3, 4'hf, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'h7, 4'hd, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h7, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0 };
assign dw_0[364] = dw_0_364[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_365 = { 4'h1, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h4, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc };
assign dw_0[365] = dw_0_365[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_366 = { 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'h7, 4'h7, 4'h1, 4'hc, 4'h3, 4'h4, 4'h0, 4'hd, 4'h4, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0 };
assign dw_0[366] = dw_0_366[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_367 = { 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'hd, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'h3, 4'h4, 4'h4, 4'hc, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h7, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[367] = dw_0_367[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_368 = { 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h4, 4'h4, 4'hf, 4'h3, 4'h3, 4'hc, 4'h3, 4'h3, 4'h1, 4'h3, 4'h0, 4'h7, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'hd, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'hf, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h1, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'hc };
assign dw_0[368] = dw_0_368[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_369 = { 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'h1, 4'h3, 4'h3, 4'hd, 4'h3, 4'hc, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h7, 4'hc, 4'h1, 4'hd, 4'h4, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc };
assign dw_0[369] = dw_0_369[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_370 = { 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'hd, 4'h1, 4'h0, 4'hc, 4'h4, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h3, 4'hd, 4'h0, 4'h7, 4'hc, 4'h0, 4'h3, 4'h0, 4'h7, 4'h3, 4'h3, 4'h0, 4'h3, 4'hd, 4'h3, 4'h3, 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc };
assign dw_0[370] = dw_0_370[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_371 = { 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'h5, 4'h7, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'h5, 4'hf, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'h7, 4'hc, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hd, 4'h1, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'hf };
assign dw_0[371] = dw_0_371[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_372 = { 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'hf, 4'h0, 4'hc, 4'hc, 4'h3, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hd, 4'hf, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'hc, 4'hd, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'hf };
assign dw_0[372] = dw_0_372[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_373 = { 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'hc, 4'h5, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hd, 4'h0, 4'h1, 4'h3, 4'h7, 4'hd, 4'h0, 4'hf, 4'hc, 4'h3, 4'h3, 4'h3, 4'hc, 4'h3, 4'hd, 4'h0, 4'hf, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'hc, 4'hf };
assign dw_0[373] = dw_0_373[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_374 = { 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h5, 4'h7, 4'hc, 4'h3, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3, 4'h0, 4'h5, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'hc, 4'h1, 4'h3, 4'h7, 4'hd, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'h1, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf };
assign dw_0[374] = dw_0_374[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_375 = { 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h7, 4'h0, 4'h1, 4'hc, 4'h0, 4'h4, 4'hf, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h3, 4'h1, 4'hf, 4'h7, 4'hd, 4'h0, 4'hf, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'hc, 4'hf, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf };
assign dw_0[375] = dw_0_375[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_376 = { 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'h1, 4'h3, 4'hc, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h1, 4'hf, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc };
assign dw_0[376] = dw_0_376[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_377 = { 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'hf, 4'h1, 4'h7, 4'hf, 4'h3, 4'hf, 4'hc, 4'h3, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h1, 4'hf, 4'h7, 4'hd, 4'h3, 4'h0, 4'h1, 4'h7, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc };
assign dw_0[377] = dw_0_377[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_378 = { 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'hf, 4'h0, 4'hc, 4'hc, 4'h3, 4'h1, 4'h0, 4'h3, 4'hc, 4'h4, 4'h0, 4'h3, 4'h3, 4'hc, 4'hc, 4'hc, 4'hc, 4'h1, 4'h3, 4'h4, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h7, 4'hc, 4'h1, 4'h5, 4'h4, 4'hf, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'hf };
assign dw_0[378] = dw_0_378[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_379 = { 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h1, 4'h3, 4'hc, 4'h1, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'hd, 4'h7, 4'h1, 4'h7, 4'h7, 4'hd, 4'h0, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h7, 4'hc, 4'h1, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'hf };
assign dw_0[379] = dw_0_379[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_380 = { 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h7, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'hc, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h7, 4'h1, 4'h0, 4'h7, 4'hc, 4'h3, 4'hf, 4'h0, 4'h7, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'hd, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'hc, 4'hf };
assign dw_0[380] = dw_0_380[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_381 = { 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hd, 4'h3, 4'h0, 4'h4, 4'hd, 4'h1, 4'h4, 4'hc, 4'hc, 4'h3, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'hf, 4'hc, 4'h1, 4'h0, 4'h3, 4'hd, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf };
assign dw_0[381] = dw_0_381[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_382 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h5, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h5, 4'hf, 4'h7, 4'hd, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf };
assign dw_0[382] = dw_0_382[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_383 = { 4'h1, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h4, 4'hc, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'hd, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h4, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h7, 4'hd, 4'h1, 4'hf, 4'h5, 4'h3, 4'h3, 4'hf, 4'hc, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'hc, 4'hd, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'hc, 4'hf };
assign dw_0[383] = dw_0_383[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_384 = { 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h3, 4'h4, 4'hf, 4'h0, 4'hc, 4'h7, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h5, 4'h1, 4'h3, 4'h4, 4'h1, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h1, 4'h7, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h5, 4'hd, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h4, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0 };
assign dw_0[384] = dw_0_384[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_385 = { 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hc, 4'h5, 4'h3, 4'h3, 4'hf, 4'h0, 4'hc, 4'h4, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'hd, 4'h3, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h1, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hf, 4'h4, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h3, 4'hd, 4'hc, 4'h5, 4'h0, 4'h0, 4'h5, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h4 };
assign dw_0[385] = dw_0_385[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_386 = { 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h5, 4'h0, 4'hc, 4'hf, 4'h3, 4'hc, 4'h4, 4'h4, 4'hc, 4'hc, 4'h3, 4'h3, 4'h5, 4'hd, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h5, 4'hd, 4'hf, 4'h0, 4'h0, 4'h1, 4'h3, 4'hf, 4'h0, 4'h4, 4'hf, 4'h3, 4'hd, 4'h3, 4'h4, 4'h0, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0 };
assign dw_0[386] = dw_0_386[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_387 = { 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'h4, 4'hc, 4'hc, 4'hf, 4'h0, 4'hc, 4'h7, 4'h1, 4'hc, 4'h0, 4'h3, 4'h3, 4'h5, 4'h1, 4'h3, 4'h4, 4'h5, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'hf, 4'h0, 4'h4, 4'h3, 4'h3, 4'hd, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0 };
assign dw_0[387] = dw_0_387[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_388 = { 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'hf, 4'h0, 4'hc, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hd, 4'h1, 4'h3, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h5, 4'h4, 4'h0, 4'hd, 4'h0, 4'h0, 4'hf, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'h0, 4'h7, 4'h0, 4'h3, 4'hd, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0 };
assign dw_0[388] = dw_0_388[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_389 = { 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'h4, 4'h4, 4'hc, 4'hc, 4'h3, 4'h3, 4'h5, 4'h1, 4'h7, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'h0, 4'hd, 4'hc, 4'hc, 4'hf, 4'h4, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h3, 4'h3, 4'hd, 4'hf, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0 };
assign dw_0[389] = dw_0_389[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_390 = { 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h5, 4'h1, 4'h3, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'hd, 4'h0, 4'h3, 4'hc, 4'hd, 4'h0, 4'hd, 4'h3, 4'h4, 4'hd, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h3, 4'h1, 4'hf, 4'h1, 4'h0, 4'h0, 4'h4, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0 };
assign dw_0[390] = dw_0_390[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_391 = { 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h4, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'hf, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'h4, 4'h5, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'hf, 4'h1, 4'h7, 4'h0, 4'hd, 4'h0, 4'h3, 4'hf, 4'h4, 4'hc, 4'hf, 4'h4, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'h7, 4'h3, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0 };
assign dw_0[391] = dw_0_391[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_392 = { 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hc, 4'h5, 4'hc, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h1, 4'h3, 4'h5, 4'h1, 4'h3, 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'hd, 4'h0, 4'h5, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h5, 4'h1, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4 };
assign dw_0[392] = dw_0_392[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_393 = { 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h4, 4'hd, 4'h0, 4'hf, 4'h0, 4'hf, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h4, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'hc, 4'h5, 4'h3, 4'hc, 4'hd, 4'h0, 4'h3, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'h3, 4'h5, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0 };
assign dw_0[393] = dw_0_393[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_394 = { 4'h3, 4'hd, 4'hc, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h4, 4'h1, 4'hc, 4'hf, 4'h0, 4'h3, 4'h1, 4'h1, 4'h3, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'hd, 4'h1, 4'h7, 4'hc, 4'hd, 4'h0, 4'h1, 4'hf, 4'h5, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'hf, 4'h4, 4'h0, 4'h0, 4'h7, 4'h7, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h4 };
assign dw_0[394] = dw_0_394[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_395 = { 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'hf, 4'h3, 4'hc, 4'h4, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'hd, 4'h1, 4'h5, 4'h0, 4'hc, 4'hd, 4'h0, 4'h0, 4'hf, 4'h5, 4'hd, 4'hf, 4'h0, 4'h1, 4'h3, 4'h0, 4'hf, 4'h0, 4'h4, 4'hc, 4'h3, 4'h5, 4'hc, 4'h1, 4'h0, 4'h3, 4'h4, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0 };
assign dw_0[395] = dw_0_395[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_396 = { 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'hf, 4'hf, 4'h3, 4'hc, 4'h4, 4'h4, 4'hc, 4'hc, 4'h0, 4'h3, 4'h1, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'hd, 4'hd, 4'h5, 4'h7, 4'h0, 4'hd, 4'h0, 4'h3, 4'hf, 4'h1, 4'hd, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'hf, 4'h0, 4'h7, 4'h0, 4'h3, 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0 };
assign dw_0[396] = dw_0_396[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_397 = { 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h1, 4'h3, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h7, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h5, 4'h1, 4'hf, 4'h0, 4'h0, 4'hd, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h3, 4'h5, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4 };
assign dw_0[397] = dw_0_397[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_398 = { 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h5, 4'h1, 4'h3, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'hd, 4'h0, 4'h3, 4'h3, 4'h4, 4'h1, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h3, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0 };
assign dw_0[398] = dw_0_398[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_399 = { 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h3, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hd, 4'h0, 4'h1, 4'hd, 4'h0, 4'hc, 4'hc, 4'h4, 4'h1, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0 };
assign dw_0[399] = dw_0_399[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_400 = { 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h7, 4'h7, 4'hc, 4'hf, 4'h3, 4'h3, 4'h5, 4'h1, 4'hd, 4'h3, 4'h1, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h4, 4'h5, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h5, 4'hc, 4'hf, 4'h7, 4'h0, 4'hd, 4'hc, 4'h7, 4'hd, 4'h1, 4'h4, 4'h5, 4'h4, 4'h3, 4'h1, 4'h0, 4'h5, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'hd, 4'h3, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc };
assign dw_0[400] = dw_0_400[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_401 = { 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h7, 4'h4, 4'hc, 4'hc, 4'h3, 4'h3, 4'h4, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h5, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h4, 4'hc, 4'hf, 4'h7, 4'h0, 4'h4, 4'hf, 4'h7, 4'h1, 4'h1, 4'h4, 4'h1, 4'h7, 4'hc, 4'h1, 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h1, 4'hd, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'h7, 4'h4, 4'hf };
assign dw_0[401] = dw_0_401[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_402 = { 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h1, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'h1, 4'hc, 4'h4, 4'hc, 4'hf, 4'h7, 4'h0, 4'h5, 4'hf, 4'h7, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'h7, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h1, 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h5, 4'h3, 4'h4, 4'hc };
assign dw_0[402] = dw_0_402[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_403 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h7, 4'hf, 4'h0, 4'h7, 4'hf, 4'h0, 4'h0, 4'hd, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'hf, 4'h3, 4'h1, 4'h0, 4'h0, 4'hd, 4'h4, 4'hf, 4'hf, 4'h4, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h1, 4'h4, 4'h1, 4'h7, 4'hc, 4'h0, 4'h0, 4'h5, 4'hd, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'h3, 4'h1, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h5, 4'h3, 4'h4, 4'hf };
assign dw_0[403] = dw_0_403[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_404 = { 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h3, 4'h7, 4'hd, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'h1, 4'hc, 4'h4, 4'hf, 4'hf, 4'h4, 4'h0, 4'h0, 4'hf, 4'h7, 4'h0, 4'h1, 4'h4, 4'h5, 4'h7, 4'h0, 4'h3, 4'h0, 4'h1, 4'hd, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h3, 4'h4, 4'hf };
assign dw_0[404] = dw_0_404[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_405 = { 4'h4, 4'hd, 4'h0, 4'h1, 4'h0, 4'h7, 4'h7, 4'hc, 4'h4, 4'h3, 4'h3, 4'h3, 4'h0, 4'hc, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h1, 4'hc, 4'hf, 4'h7, 4'h0, 4'h0, 4'hf, 4'h7, 4'hc, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h1, 4'hd, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf };
assign dw_0[405] = dw_0_405[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_406 = { 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h7, 4'h7, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'hc, 4'hf, 4'h7, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'h5, 4'hf, 4'h1, 4'h0, 4'h5, 4'hd, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'hf, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0 };
assign dw_0[406] = dw_0_406[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_407 = { 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'hd, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h4, 4'h3, 4'h1, 4'h5, 4'h1, 4'h5, 4'h4, 4'h0, 4'h3, 4'hc, 4'h1, 4'h4, 4'hd, 4'hc, 4'h4, 4'hf, 4'hf, 4'h7, 4'h0, 4'h0, 4'hf, 4'h7, 4'h1, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'h3, 4'h5, 4'h3, 4'h0, 4'h0, 4'h3, 4'h1, 4'h5, 4'hf, 4'hc, 4'h0, 4'h0, 4'h5, 4'h3, 4'h4, 4'hc };
assign dw_0[407] = dw_0_407[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_408 = { 4'h7, 4'hc, 4'hc, 4'h1, 4'h0, 4'h7, 4'h4, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'h1, 4'hd, 4'h3, 4'hc, 4'h3, 4'h3, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'h4, 4'hf, 4'hc, 4'h0, 4'h4, 4'h0, 4'hd, 4'h4, 4'hf, 4'hf, 4'h7, 4'h0, 4'h1, 4'hf, 4'h3, 4'hc, 4'h1, 4'h4, 4'h1, 4'h7, 4'hc, 4'hc, 4'h0, 4'h5, 4'hc, 4'h3, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'hd, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'hf };
assign dw_0[408] = dw_0_408[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_409 = { 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h7, 4'h4, 4'hc, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'hd, 4'h3, 4'hc, 4'h0, 4'h3, 4'h1, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'hd, 4'h4, 4'hc, 4'hf, 4'h7, 4'h4, 4'h0, 4'hf, 4'h7, 4'hc, 4'h1, 4'h4, 4'h1, 4'h4, 4'hf, 4'h0, 4'h0, 4'h5, 4'hc, 4'h3, 4'hd, 4'h7, 4'h5, 4'hc, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc };
assign dw_0[409] = dw_0_409[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_410 = { 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'hf, 4'h4, 4'h3, 4'hc, 4'h0, 4'h1, 4'hd, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h1, 4'h1, 4'h4, 4'h5, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'hf, 4'hf, 4'h4, 4'h3, 4'h1, 4'hf, 4'h7, 4'hc, 4'h1, 4'h0, 4'h1, 4'h5, 4'hf, 4'h0, 4'h0, 4'h5, 4'hd, 4'h0, 4'hd, 4'h3, 4'h4, 4'h0, 4'h3, 4'h1, 4'h1, 4'hf, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'h4, 4'hc };
assign dw_0[410] = dw_0_410[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_411 = { 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'h3, 4'h4, 4'hc, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'hd, 4'hf, 4'h1, 4'h0, 4'h0, 4'h1, 4'h5, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h4, 4'hc, 4'hf, 4'h7, 4'h0, 4'h1, 4'hf, 4'h4, 4'h0, 4'hc, 4'h4, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'hd, 4'h0, 4'hc, 4'h7, 4'h1, 4'h0, 4'h7, 4'h1, 4'h5, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'h4, 4'hc };
assign dw_0[411] = dw_0_411[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_412 = { 4'h4, 4'hc, 4'h0, 4'h1, 4'h0, 4'h7, 4'h4, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h4, 4'h5, 4'h4, 4'h3, 4'h3, 4'hd, 4'h0, 4'h0, 4'hc, 4'h4, 4'hf, 4'hf, 4'h7, 4'h0, 4'h0, 4'hf, 4'h7, 4'h4, 4'hd, 4'h4, 4'h5, 4'h4, 4'hc, 4'h1, 4'h0, 4'h1, 4'hd, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'hd, 4'h5, 4'h7, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'hf };
assign dw_0[412] = dw_0_412[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_413 = { 4'h5, 4'hd, 4'h0, 4'h1, 4'h0, 4'h7, 4'h4, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h5, 4'h1, 4'h4, 4'h5, 4'h0, 4'h3, 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'hf, 4'h7, 4'h0, 4'h0, 4'hf, 4'h4, 4'h4, 4'h1, 4'h0, 4'h1, 4'h4, 4'hc, 4'h1, 4'h0, 4'h1, 4'hc, 4'h7, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h3, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'hc };
assign dw_0[413] = dw_0_413[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_414 = { 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h7, 4'hd, 4'hc, 4'h3, 4'h3, 4'h4, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h4, 4'h4, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hd, 4'h4, 4'hc, 4'hf, 4'h7, 4'h0, 4'h5, 4'hc, 4'h4, 4'h0, 4'h1, 4'h4, 4'h1, 4'h7, 4'h1, 4'h1, 4'h0, 4'h5, 4'hd, 4'h3, 4'hc, 4'h3, 4'h1, 4'h0, 4'h3, 4'h1, 4'h5, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'hf };
assign dw_0[414] = dw_0_414[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_415 = { 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'h3, 4'h7, 4'hd, 4'hc, 4'h3, 4'h3, 4'h0, 4'hf, 4'hd, 4'h3, 4'hd, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h5, 4'hd, 4'h4, 4'hc, 4'hf, 4'h7, 4'h0, 4'h5, 4'hf, 4'h4, 4'h5, 4'h0, 4'h4, 4'h5, 4'h7, 4'hc, 4'hc, 4'h0, 4'h1, 4'hc, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h7, 4'h4, 4'hf };
assign dw_0[415] = dw_0_415[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_416 = { 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h5, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h3, 4'h3, 4'h3, 4'hf, 4'h5, 4'hc, 4'h4, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'h7, 4'h7, 4'h1, 4'h5, 4'h5, 4'h1, 4'h0, 4'hc, 4'hc, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hc, 4'h3, 4'hc, 4'hc, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'h7, 4'h1, 4'h0, 4'h3, 4'hc, 4'hc, 4'h4 };
assign dw_0[416] = dw_0_416[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_417 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h1, 4'h1, 4'h0, 4'h0, 4'h3, 4'h7, 4'hc, 4'h4, 4'h5, 4'h1, 4'h0, 4'h1, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h4, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0 };
assign dw_0[417] = dw_0_417[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_418 = { 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'hd, 4'hd, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h7, 4'h3, 4'h7, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h4, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'hf, 4'hc, 4'hc, 4'hf, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0 };
assign dw_0[418] = dw_0_418[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_419 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h3, 4'hc, 4'h0, 4'hd, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'h4, 4'h5, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'hf, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0 };
assign dw_0[419] = dw_0_419[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_420 = { 4'h0, 4'h7, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h7, 4'h4, 4'hc, 4'h0, 4'hc, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h4, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[420] = dw_0_420[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_421 = { 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h4, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'hf, 4'h1, 4'h4, 4'h0, 4'h3, 4'h3, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[421] = dw_0_421[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_422 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hd, 4'h4, 4'h0, 4'h3, 4'h1, 4'hc, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h1, 4'hc, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[422] = dw_0_422[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_423 = { 4'hc, 4'h7, 4'h4, 4'h1, 4'h0, 4'h1, 4'h4, 4'h7, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h4, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h7, 4'hc, 4'h7, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[423] = dw_0_423[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_424 = { 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h7, 4'h1, 4'h7, 4'h5, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0 };
assign dw_0[424] = dw_0_424[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_425 = { 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h4, 4'hc, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h7, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0 };
assign dw_0[425] = dw_0_425[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_426 = { 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h7, 4'h0, 4'hc, 4'h3, 4'hc, 4'h4, 4'h4, 4'h1, 4'h3, 4'h0, 4'h0, 4'h7, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'hc, 4'h0, 4'h0, 4'hc, 4'h4, 4'h3, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'hd, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h1, 4'h7, 4'h0, 4'h3, 4'hf, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7 };
assign dw_0[426] = dw_0_426[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_427 = { 4'hc, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'h4, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0 };
assign dw_0[427] = dw_0_427[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_428 = { 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'hc, 4'hc, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0 };
assign dw_0[428] = dw_0_428[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_429 = { 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'hc, 4'h4, 4'h5, 4'h1, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h1, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4 };
assign dw_0[429] = dw_0_429[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_430 = { 4'hc, 4'h7, 4'h0, 4'h1, 4'h0, 4'h1, 4'hd, 4'h7, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h4, 4'h0, 4'h4, 4'hc, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'hf, 4'hf, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h3, 4'h3, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0 };
assign dw_0[430] = dw_0_430[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_431 = { 4'hc, 4'h4, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'hf, 4'h0, 4'hc, 4'hc, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'h5, 4'h5, 4'hd, 4'h0, 4'h3, 4'h0, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'hf, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0 };
assign dw_0[431] = dw_0_431[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_432 = { 4'h0, 4'hd, 4'h4, 4'h1, 4'h0, 4'h1, 4'h4, 4'h5, 4'hc, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h7, 4'h5, 4'hf, 4'h3, 4'hd, 4'h0, 4'h7, 4'h4, 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc, 4'hf, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h1, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'hd, 4'h1, 4'hc, 4'h0, 4'h0, 4'h7, 4'h5, 4'h0, 4'h7, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h1 };
assign dw_0[432] = dw_0_432[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_433 = { 4'h0, 4'hd, 4'h4, 4'h1, 4'h0, 4'hd, 4'h3, 4'h5, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h7, 4'h4, 4'hc, 4'h0, 4'hd, 4'h1, 4'h4, 4'h4, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'hd, 4'h0, 4'hc, 4'hf, 4'hc, 4'h3, 4'h0, 4'hc, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h7, 4'h0, 4'h3, 4'hd, 4'h1, 4'hf, 4'h0, 4'h0, 4'h7, 4'h5, 4'h3, 4'h3, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h4 };
assign dw_0[433] = dw_0_433[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_434 = { 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'h3, 4'h4, 4'hd, 4'h0, 4'hd, 4'h1, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h1, 4'hc, 4'h0, 4'hd, 4'hd, 4'hf, 4'hc, 4'hf, 4'h0, 4'h3, 4'h3, 4'hc, 4'h5, 4'h0, 4'h4, 4'hc, 4'h0, 4'h1, 4'hd, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hd, 4'hd, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4 };
assign dw_0[434] = dw_0_434[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_435 = { 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'hc, 4'h0, 4'h1, 4'hd, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'h3, 4'hc, 4'h4, 4'h7, 4'h0, 4'hc, 4'h0, 4'h1, 4'hd, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'hf, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h5, 4'h0, 4'hc, 4'h4 };
assign dw_0[435] = dw_0_435[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_436 = { 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'h3, 4'h4, 4'h4, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'hd, 4'h0, 4'hc, 4'hf, 4'hc, 4'h0, 4'hc, 4'hc, 4'h1, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'hd, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'hd, 4'h1, 4'hc, 4'h0, 4'h0, 4'h7, 4'h5, 4'h3, 4'h3, 4'h1, 4'h0, 4'h7, 4'h0, 4'h4, 4'h0 };
assign dw_0[436] = dw_0_436[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_437 = { 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'h4, 4'h3, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'h4, 4'h0, 4'h3, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h1, 4'h0, 4'h4, 4'h1, 4'hd, 4'hc, 4'hd, 4'hf, 4'hc, 4'h1, 4'hf, 4'hc, 4'h5, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'h0, 4'h7, 4'h4, 4'h7, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h3 };
assign dw_0[437] = dw_0_437[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_438 = { 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'h1, 4'h3, 4'hd, 4'h5, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'hd, 4'h0, 4'h3, 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'hd, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h1, 4'hd, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h1, 4'hc, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h3 };
assign dw_0[438] = dw_0_438[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_439 = { 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h4, 4'h7, 4'h1, 4'h4, 4'h0, 4'hd, 4'h3, 4'h0, 4'h7, 4'h3, 4'h4, 4'h1, 4'h1, 4'hd, 4'h0, 4'h3, 4'h0, 4'h7, 4'h4, 4'h1, 4'h1, 4'h0, 4'h4, 4'h1, 4'hd, 4'h3, 4'h0, 4'hf, 4'hc, 4'h1, 4'h3, 4'hc, 4'h4, 4'h0, 4'hc, 4'hc, 4'hf, 4'h3, 4'hd, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h5, 4'hd, 4'hc, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc, 4'hc, 4'h3 };
assign dw_0[439] = dw_0_439[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_440 = { 4'hc, 4'hd, 4'h0, 4'h1, 4'h0, 4'h1, 4'h7, 4'h5, 4'h4, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h1, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'h4, 4'h4, 4'h1, 4'h1, 4'hc, 4'h4, 4'h1, 4'hd, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'h4, 4'h3, 4'hd, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h5, 4'h1, 4'hf, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3 };
assign dw_0[440] = dw_0_440[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_441 = { 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h1, 4'h7, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h7, 4'h3, 4'h4, 4'h1, 4'h3, 4'hd, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'hd, 4'h1, 4'h0, 4'h4, 4'h1, 4'hd, 4'hc, 4'hc, 4'hf, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h4, 4'h3, 4'hd, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'h5, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[441] = dw_0_441[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_442 = { 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'h0, 4'h7, 4'h5, 4'h4, 4'h1, 4'h1, 4'h3, 4'hc, 4'h4, 4'h3, 4'h4, 4'h1, 4'h3, 4'hc, 4'h1, 4'h3, 4'h4, 4'h7, 4'h4, 4'h1, 4'h1, 4'hc, 4'h4, 4'h1, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'h1, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h5, 4'h1, 4'hf, 4'h0, 4'h0, 4'h7, 4'h4, 4'h7, 4'h0, 4'h1, 4'h0, 4'h7, 4'hc, 4'hc, 4'h3 };
assign dw_0[442] = dw_0_442[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_443 = { 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h1, 4'h1, 4'hc, 4'h4, 4'hd, 4'hd, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h1, 4'hc, 4'h0, 4'h4, 4'h7, 4'h4, 4'h3, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'hc, 4'h0 };
assign dw_0[443] = dw_0_443[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_444 = { 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'hc, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'hd, 4'hd, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h1, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h1, 4'hc, 4'h0, 4'h0, 4'h7, 4'h4, 4'h7, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3 };
assign dw_0[444] = dw_0_444[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_445 = { 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h0, 4'h4, 4'h4, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'hd, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h7, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hd, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h5, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0 };
assign dw_0[445] = dw_0_445[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_446 = { 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h7, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'hd, 4'hc, 4'h0, 4'hc, 4'hf, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h1, 4'hd, 4'h0, 4'h3, 4'h7, 4'h5, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'h5 };
assign dw_0[446] = dw_0_446[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_447 = { 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'h1, 4'h7, 4'h1, 4'h3, 4'hd, 4'h4, 4'h0, 4'hc, 4'h3, 4'h7, 4'h4, 4'hc, 4'h3, 4'hd, 4'h4, 4'h3, 4'h0, 4'h7, 4'h4, 4'h1, 4'h5, 4'hc, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc, 4'hf, 4'hd, 4'h3, 4'hf, 4'hd, 4'h4, 4'hc, 4'h4, 4'hc, 4'h4, 4'h1, 4'hd, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'h1, 4'hc, 4'h0, 4'h3, 4'h3, 4'h5, 4'h3, 4'h7, 4'h5, 4'h0, 4'h7, 4'hc, 4'h0, 4'h1 };
assign dw_0[447] = dw_0_447[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_448 = { 4'hd, 4'h7, 4'hc, 4'h0, 4'h0, 4'hd, 4'hd, 4'h7, 4'h4, 4'h1, 4'hc, 4'h5, 4'h7, 4'h0, 4'h4, 4'h7, 4'h1, 4'h1, 4'h3, 4'h1, 4'hc, 4'hf, 4'h1, 4'hc, 4'hc, 4'h3, 4'hc, 4'h4, 4'h3, 4'h4, 4'h5, 4'h3, 4'h4, 4'h1, 4'hc, 4'h4, 4'hf, 4'h7, 4'h3, 4'hf, 4'h0, 4'hc, 4'h7, 4'hd, 4'h3, 4'h3, 4'h3, 4'hd, 4'h0, 4'hf, 4'h5, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf };
assign dw_0[448] = dw_0_448[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_449 = { 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h7, 4'h3, 4'h1, 4'hd, 4'h5, 4'h7, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'h4, 4'h4, 4'hd, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h1, 4'h3, 4'h7, 4'hd, 4'h3, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'hd, 4'h3, 4'h0, 4'hc, 4'hd, 4'h0, 4'h3, 4'h1, 4'hf, 4'h0, 4'h3, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'hc, 4'hf };
assign dw_0[449] = dw_0_449[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_450 = { 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h3, 4'h1, 4'hc, 4'h4, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h3, 4'h7, 4'hd, 4'h3, 4'hf, 4'hf, 4'h7, 4'h3, 4'h1, 4'h0, 4'h3, 4'h3, 4'hc, 4'h7, 4'h3, 4'h3, 4'hd, 4'h0, 4'h3, 4'h5, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'hf };
assign dw_0[450] = dw_0_450[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_451 = { 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h7, 4'h3, 4'h1, 4'hd, 4'h0, 4'h4, 4'h3, 4'h4, 4'h4, 4'h3, 4'h0, 4'h1, 4'h0, 4'hd, 4'hc, 4'h4, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'hd, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'hd, 4'h3, 4'h3, 4'h3, 4'hd, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0 };
assign dw_0[451] = dw_0_451[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_452 = { 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h7, 4'h3, 4'h1, 4'h0, 4'h1, 4'h4, 4'h3, 4'h4, 4'h4, 4'h3, 4'h0, 4'h3, 4'h3, 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h7, 4'h1, 4'h3, 4'h4, 4'hd, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'hd, 4'h4, 4'h0, 4'h3, 4'hd, 4'h3, 4'hc, 4'h1, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'hc };
assign dw_0[452] = dw_0_452[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_453 = { 4'h1, 4'h7, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h7, 4'h3, 4'h1, 4'hd, 4'h5, 4'h4, 4'h3, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h1, 4'h3, 4'h4, 4'hd, 4'h3, 4'h3, 4'hc, 4'h7, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'h7, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'hc };
assign dw_0[453] = dw_0_453[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_454 = { 4'h1, 4'h7, 4'hc, 4'h0, 4'h0, 4'h1, 4'hd, 4'h4, 4'h3, 4'h1, 4'h1, 4'h5, 4'h4, 4'h3, 4'h4, 4'h4, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h7, 4'hd, 4'h3, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'hf, 4'h5, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc };
assign dw_0[454] = dw_0_454[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_455 = { 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h1, 4'h1, 4'h5, 4'h4, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'hd, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h5, 4'hc, 4'h0, 4'h3, 4'hf, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[455] = dw_0_455[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_456 = { 4'h1, 4'h7, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h3, 4'hd, 4'hd, 4'h5, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h1, 4'h3, 4'h7, 4'h1, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hd, 4'h0, 4'hf, 4'h5, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h7, 4'h1, 4'h0, 4'h3, 4'h1, 4'hc, 4'hf };
assign dw_0[456] = dw_0_456[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_457 = { 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h7, 4'h3, 4'h0, 4'h1, 4'h4, 4'h4, 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h1, 4'h3, 4'h0, 4'hc, 4'h3, 4'hc, 4'h4, 4'h0, 4'h3, 4'hf, 4'hd, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'hc, 4'h1, 4'hf, 4'h0, 4'h3, 4'h3, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h1, 4'hc, 4'hf };
assign dw_0[457] = dw_0_457[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_458 = { 4'hc, 4'h7, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h7, 4'hf, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h1, 4'h3, 4'h7, 4'hd, 4'h0, 4'h3, 4'hc, 4'hc, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3 };
assign dw_0[458] = dw_0_458[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_459 = { 4'h1, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'h1, 4'h1, 4'h1, 4'h4, 4'h3, 4'h4, 4'h4, 4'h3, 4'h0, 4'h4, 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h7, 4'h1, 4'h3, 4'h7, 4'hd, 4'h3, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h3, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h5, 4'hf, 4'h0, 4'h3, 4'hf, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h3 };
assign dw_0[459] = dw_0_459[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_460 = { 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h1, 4'h7, 4'h3, 4'h1, 4'hd, 4'h4, 4'h4, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h3, 4'h7, 4'h1, 4'h3, 4'hc, 4'hf, 4'h3, 4'hc, 4'h0, 4'hc, 4'h3, 4'h3, 4'hd, 4'h0, 4'h0, 4'h7, 4'hc, 4'h0, 4'hf, 4'h1, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'h4, 4'h3, 4'h1, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3 };
assign dw_0[460] = dw_0_460[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_461 = { 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'hd, 4'hd, 4'h7, 4'h3, 4'h1, 4'h1, 4'h1, 4'h4, 4'h4, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'hd, 4'hc, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h7, 4'hd, 4'h3, 4'h3, 4'hf, 4'h4, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'hf, 4'hd, 4'h0, 4'hf, 4'h5, 4'hf, 4'h0, 4'h3, 4'h3, 4'h1, 4'h4, 4'h7, 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0 };
assign dw_0[461] = dw_0_461[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_462 = { 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'h7, 4'h1, 4'h1, 4'h5, 4'h4, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'hd, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'h0, 4'h3, 4'hd, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc, 4'h3, 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h7, 4'h1, 4'hc, 4'h0 };
assign dw_0[462] = dw_0_462[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_463 = { 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h7, 4'h3, 4'h1, 4'hc, 4'h0, 4'h4, 4'h3, 4'h4, 4'h4, 4'hc, 4'h0, 4'h7, 4'h3, 4'hd, 4'hc, 4'h4, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h1, 4'h0, 4'h7, 4'hd, 4'h0, 4'h3, 4'hf, 4'h0, 4'hc, 4'hc, 4'hc, 4'hf, 4'h3, 4'hc, 4'h3, 4'h3, 4'hf, 4'hc, 4'h3, 4'hf, 4'h1, 4'h3, 4'h0, 4'h3, 4'hf, 4'hc, 4'h4, 4'h4, 4'h5, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0 };
assign dw_0[463] = dw_0_463[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_464 = { 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h3, 4'hf, 4'h5, 4'hc, 4'h4, 4'h0, 4'hd, 4'h7, 4'h4, 4'h3, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h5, 4'h3, 4'h4, 4'h0, 4'h7, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'h1, 4'h1, 4'hc, 4'hf };
assign dw_0[464] = dw_0_464[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_465 = { 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'hf, 4'h4, 4'h0, 4'h5, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'hd, 4'h3, 4'h0, 4'hc, 4'h1, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h5, 4'h3, 4'h0, 4'hc, 4'h3, 4'hd, 4'h0, 4'h3, 4'hc, 4'h7, 4'h3, 4'h3, 4'h4, 4'h0, 4'h1, 4'hf, 4'h7, 4'h0, 4'h7, 4'h1, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'hc, 4'hf };
assign dw_0[465] = dw_0_465[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_466 = { 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h4, 4'hc, 4'h5, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h7, 4'hd, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'h4, 4'h4, 4'h3, 4'h0, 4'h3, 4'h7, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf };
assign dw_0[466] = dw_0_466[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_467 = { 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h4, 4'h5, 4'h1, 4'h5, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'h4, 4'hf, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h7, 4'h0, 4'h3, 4'hd, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf };
assign dw_0[467] = dw_0_467[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_468 = { 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'hc, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'hc, 4'h3, 4'hd, 4'h0, 4'hf, 4'hc, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'h1, 4'h7, 4'h3, 4'h0, 4'h0, 4'h5, 4'h1, 4'hc, 4'hc };
assign dw_0[468] = dw_0_468[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_469 = { 4'h1, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h5, 4'h0, 4'h5, 4'h4, 4'hc, 4'h7, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h3, 4'h3, 4'h1, 4'h0, 4'h1, 4'hc, 4'h4, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'hc, 4'hc };
assign dw_0[469] = dw_0_469[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_470 = { 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h4, 4'hd, 4'h5, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'hc, 4'hd, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h7, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf };
assign dw_0[470] = dw_0_470[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_471 = { 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h5, 4'hc, 4'h4, 4'h4, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h4, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'h0, 4'h4, 4'h1, 4'h1, 4'hf, 4'h7, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h4, 4'hd, 4'h0, 4'h3, 4'h4, 4'h4, 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc };
assign dw_0[471] = dw_0_471[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_472 = { 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h4, 4'hd, 4'h5, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'hf, 4'h7, 4'h3, 4'h3, 4'h4, 4'h1, 4'h0, 4'hc, 4'h7, 4'h0, 4'h3, 4'h5, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf };
assign dw_0[472] = dw_0_472[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_473 = { 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h5, 4'hc, 4'h5, 4'h0, 4'hc, 4'h4, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc, 4'h0, 4'hd, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h7, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h7, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'hf };
assign dw_0[473] = dw_0_473[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_474 = { 4'h1, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h5, 4'hd, 4'h5, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h1, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc, 4'h3, 4'hc, 4'h3, 4'hf, 4'hc, 4'h7, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hf, 4'h7, 4'h0, 4'h3, 4'h1, 4'h1, 4'h5, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'hf };
assign dw_0[474] = dw_0_474[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_475 = { 4'h1, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h5, 4'hd, 4'h5, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'hc, 4'hd, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'hd, 4'h0, 4'h3, 4'hc, 4'h3, 4'h7, 4'h3, 4'h4, 4'h0, 4'h0, 4'hf, 4'h7, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3, 4'h4, 4'hd, 4'h0, 4'h0, 4'h7, 4'h5, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf };
assign dw_0[475] = dw_0_475[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_476 = { 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h4, 4'hd, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'hf, 4'h7, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'hf, 4'h7, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'hc, 4'hc };
assign dw_0[476] = dw_0_476[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_477 = { 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h3, 4'h4, 4'h5, 4'h1, 4'h5, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hd, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h7, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'hf };
assign dw_0[477] = dw_0_477[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_478 = { 4'h1, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h5, 4'hd, 4'h5, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h3, 4'hd, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'h3, 4'h4, 4'h7, 4'h0, 4'hf, 4'h7, 4'h0, 4'h7, 4'h1, 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf };
assign dw_0[478] = dw_0_478[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_479 = { 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'h4, 4'h5, 4'hd, 4'h4, 4'hd, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'hf, 4'h7, 4'h4, 4'h0, 4'h5, 4'h1, 4'h4, 4'hc, 4'hf, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'hf, 4'h7, 4'h1, 4'h3, 4'h5, 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0, 4'h4, 4'h4, 4'h0, 4'h5, 4'h1, 4'hc, 4'hc };
assign dw_0[479] = dw_0_479[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_480 = { 4'h7, 4'hd, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h3, 4'hf, 4'h4, 4'h1, 4'hc, 4'h1, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'hc, 4'h5, 4'h1, 4'hf, 4'h0, 4'hc, 4'h3, 4'h7, 4'h0, 4'hc, 4'h5, 4'h3, 4'h3, 4'hc, 4'hd, 4'hf, 4'h5, 4'h0, 4'h0, 4'hd, 4'hc, 4'hc, 4'h1, 4'h5, 4'h4, 4'h4, 4'h1, 4'h0, 4'h5, 4'h4, 4'h1, 4'hc, 4'h4, 4'hc, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1 };
assign dw_0[480] = dw_0_480[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_481 = { 4'h4, 4'hd, 4'h0, 4'h1, 4'h0, 4'h7, 4'h7, 4'hd, 4'h0, 4'hc, 4'h4, 4'h1, 4'hd, 4'h1, 4'h5, 4'h0, 4'h3, 4'h3, 4'hc, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'h0, 4'hd, 4'h5, 4'h3, 4'h3, 4'hc, 4'hd, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'hf, 4'hc, 4'h1, 4'h1, 4'h1, 4'h0, 4'h1, 4'h1, 4'h5, 4'h0, 4'hc, 4'h0, 4'h5, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1 };
assign dw_0[481] = dw_0_481[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_482 = { 4'h4, 4'hd, 4'h0, 4'h1, 4'h0, 4'h7, 4'h3, 4'h0, 4'h4, 4'hd, 4'h4, 4'h1, 4'hd, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'hc, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h5, 4'h3, 4'h7, 4'hd, 4'hd, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'h1, 4'h1, 4'h1, 4'h3, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h7, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1 };
assign dw_0[482] = dw_0_482[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_483 = { 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'hc, 4'h5, 4'h0, 4'h3, 4'h0, 4'hd, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'hc, 4'h0, 4'h7, 4'h3, 4'h0, 4'h5, 4'h0, 4'h7, 4'h1, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'hc, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h3, 4'h5, 4'h1, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5 };
assign dw_0[483] = dw_0_483[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_484 = { 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h7, 4'hd, 4'h1, 4'hc, 4'hf, 4'h1, 4'hd, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h5, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h7, 4'hd, 4'h5, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[484] = dw_0_484[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_485 = { 4'h7, 4'hd, 4'h0, 4'h1, 4'h0, 4'h7, 4'h7, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'hd, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hd, 4'h4, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h1, 4'h5, 4'hd, 4'hc, 4'h0, 4'hc, 4'h7, 4'h1, 4'h0, 4'h1, 4'h5, 4'h4, 4'h1, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h7, 4'h5, 4'hd, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[485] = dw_0_485[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_486 = { 4'h7, 4'hd, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'hc, 4'hd, 4'h1, 4'hf, 4'h1, 4'hd, 4'hd, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hf, 4'h5, 4'h4, 4'hc, 4'hd, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h5, 4'h1, 4'h3, 4'h0, 4'h1, 4'hd, 4'hf, 4'h0, 4'hc, 4'h7, 4'hc, 4'h0, 4'h1, 4'h1, 4'h4, 4'h1, 4'h4, 4'h0, 4'h5, 4'h0, 4'h1, 4'h7, 4'h5, 4'hd, 4'h5, 4'h4, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0 };
assign dw_0[486] = dw_0_486[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_487 = { 4'h7, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'hd, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h7, 4'h0, 4'h0, 4'h4, 4'h1, 4'h3, 4'h0, 4'h1, 4'h1, 4'hf, 4'h0, 4'hc, 4'h7, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h1, 4'h5, 4'h0, 4'h5, 4'h4, 4'h1, 4'h4, 4'h5, 4'h1, 4'h5, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[487] = dw_0_487[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_488 = { 4'h7, 4'h1, 4'hc, 4'h0, 4'h0, 4'h7, 4'h7, 4'hc, 4'h1, 4'h0, 4'hf, 4'h1, 4'hd, 4'h1, 4'h1, 4'h4, 4'h1, 4'h1, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h7, 4'h0, 4'h0, 4'h5, 4'h1, 4'h3, 4'h0, 4'h1, 4'h1, 4'hf, 4'h0, 4'hd, 4'h7, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h1, 4'h5, 4'h0, 4'h5, 4'h4, 4'h0, 4'h7, 4'h5, 4'h0, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[488] = dw_0_488[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_489 = { 4'h7, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h1, 4'h0, 4'hf, 4'h0, 4'hd, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h4, 4'hc, 4'h1, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h7, 4'h0, 4'h0, 4'h5, 4'h1, 4'h3, 4'h1, 4'h1, 4'h1, 4'h3, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h1, 4'h4, 4'h5, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h5, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0 };
assign dw_0[489] = dw_0_489[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_490 = { 4'h4, 4'hd, 4'hc, 4'h0, 4'h0, 4'h4, 4'h7, 4'hd, 4'h0, 4'hc, 4'hc, 4'h1, 4'hd, 4'h1, 4'h5, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h3, 4'h0, 4'h1, 4'hd, 4'hc, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h4, 4'h5, 4'h0, 4'h5, 4'h4, 4'h1, 4'h7, 4'h5, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[490] = dw_0_490[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_491 = { 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h1, 4'hc, 4'hd, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'hc, 4'h7, 4'h3, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'hd, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h7, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h1, 4'h3, 4'h5, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[491] = dw_0_491[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_492 = { 4'h4, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'h1, 4'h0, 4'h5, 4'hd, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'hc, 4'h3, 4'h7, 4'h0, 4'hd, 4'h1, 4'h0, 4'h7, 4'hd, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'h5, 4'hc, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1 };
assign dw_0[492] = dw_0_492[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_493 = { 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'hc, 4'h4, 4'h0, 4'h4, 4'h4, 4'hd, 4'h1, 4'h5, 4'h3, 4'h7, 4'h1, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'hf, 4'h7, 4'h3, 4'h0, 4'h1, 4'h5, 4'h3, 4'h4, 4'hc, 4'hd, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'h3, 4'h4, 4'h1, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1 };
assign dw_0[493] = dw_0_493[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_494 = { 4'h4, 4'hd, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h1, 4'h4, 4'h1, 4'h4, 4'h5, 4'hd, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h4, 4'h4, 4'h0, 4'h4, 4'hd, 4'h3, 4'h3, 4'h0, 4'h1, 4'h5, 4'h3, 4'h3, 4'hc, 4'hd, 4'hc, 4'h4, 4'h0, 4'h1, 4'h1, 4'h3, 4'h7, 4'h1, 4'h1, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h7, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1 };
assign dw_0[494] = dw_0_494[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_495 = { 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'hd, 4'h5, 4'h0, 4'h4, 4'h1, 4'hd, 4'h1, 4'h5, 4'hf, 4'h0, 4'h3, 4'h0, 4'h1, 4'h5, 4'h4, 4'hc, 4'h0, 4'h5, 4'h4, 4'hc, 4'h4, 4'hc, 4'h3, 4'h3, 4'h0, 4'hc, 4'h5, 4'h3, 4'h0, 4'hc, 4'hd, 4'hc, 4'h7, 4'h0, 4'h5, 4'hd, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h1, 4'h1, 4'h5, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd };
assign dw_0[495] = dw_0_495[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_496 = { 4'h0, 4'hd, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'hd, 4'hc, 4'hd, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'h4, 4'h5, 4'h0, 4'h7, 4'hc, 4'h4, 4'h0, 4'hd, 4'h3, 4'h4, 4'h0 };
assign dw_0[496] = dw_0_496[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_497 = { 4'h0, 4'h5, 4'hc, 4'h3, 4'h0, 4'h3, 4'h1, 4'hc, 4'hf, 4'h3, 4'h0, 4'h3, 4'h7, 4'hc, 4'h0, 4'h4, 4'h3, 4'h3, 4'h4, 4'h3, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h4, 4'hc, 4'h4, 4'h4, 4'h0, 4'h1, 4'hd, 4'h4, 4'h3, 4'hd, 4'h3, 4'h3, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h1, 4'h0, 4'h5, 4'hc, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'h1, 4'h3, 4'h4, 4'hc, 4'h0, 4'h0, 4'hd, 4'h3, 4'h4, 4'hc };
assign dw_0[497] = dw_0_497[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_498 = { 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h3, 4'h1, 4'hc, 4'h4, 4'hd, 4'h3, 4'h3, 4'h0, 4'h0, 4'h5, 4'h3, 4'hc, 4'h0, 4'hc, 4'h4, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h4, 4'h3, 4'h1, 4'h0, 4'hf, 4'h0, 4'h1, 4'hc, 4'h1, 4'h4, 4'h3, 4'h1, 4'h3, 4'h5, 4'hf, 4'h3, 4'h3, 4'h3, 4'h1, 4'h0, 4'h3, 4'h1, 4'h3, 4'h7, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'hc };
assign dw_0[498] = dw_0_498[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_499 = { 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h3, 4'hd, 4'h4, 4'hd, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0, 4'h1, 4'h3, 4'h0, 4'hc, 4'hd, 4'h4, 4'h0, 4'hd, 4'h0, 4'h3, 4'h1, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'h5, 4'h3, 4'h5, 4'h0, 4'h3, 4'h0, 4'h3, 4'h5, 4'h0, 4'h3, 4'h5, 4'hf, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'hc };
assign dw_0[499] = dw_0_499[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_500 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'h3, 4'h3, 4'h3, 4'hf, 4'h4, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h1, 4'h4, 4'hc, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'hd, 4'h4, 4'h3, 4'hc, 4'h0, 4'hf, 4'h5, 4'h1, 4'h0, 4'h1, 4'h7, 4'h3, 4'h1, 4'h3, 4'h5, 4'h3, 4'h3, 4'h3, 4'hf, 4'h1, 4'h0, 4'h0, 4'h5, 4'h7, 4'h7, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'hc };
assign dw_0[500] = dw_0_500[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_501 = { 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'hd, 4'hc, 4'h3, 4'h3, 4'h0, 4'hc, 4'h7, 4'hc, 4'hf, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hd, 4'h4, 4'hc, 4'h0, 4'h7, 4'hf, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'hd, 4'h4, 4'h3, 4'hd, 4'h0, 4'h3, 4'h5, 4'h1, 4'h4, 4'h1, 4'h4, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h5, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'h3, 4'h4, 4'hc };
assign dw_0[501] = dw_0_501[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_502 = { 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h7, 4'hc, 4'hd, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h4, 4'h3, 4'hc, 4'h0, 4'hf, 4'h1, 4'h1, 4'h0, 4'h5, 4'h4, 4'h3, 4'h1, 4'h0, 4'h5, 4'h0, 4'h3, 4'h3, 4'h3, 4'h1, 4'h0, 4'h0, 4'h5, 4'h3, 4'h7, 4'hf, 4'h0, 4'h0, 4'hd, 4'h3, 4'h4, 4'hc };
assign dw_0[502] = dw_0_502[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_503 = { 4'h0, 4'hd, 4'h4, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'h3, 4'hf, 4'h7, 4'hf, 4'h4, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'hd, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h1, 4'hc, 4'h5, 4'h0, 4'h1, 4'h3, 4'hf, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h3, 4'h1, 4'h0, 4'h5, 4'h0, 4'h7, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h5, 4'h7, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'h3, 4'h4, 4'hc };
assign dw_0[503] = dw_0_503[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_504 = { 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'hf, 4'h7, 4'hf, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'hd, 4'h4, 4'h7, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'hc, 4'h4, 4'h3, 4'hc, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'hc, 4'hd, 4'h0, 4'h5, 4'h0, 4'h3, 4'h7, 4'h3, 4'h1, 4'h0, 4'h0, 4'h5, 4'h3, 4'h4, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'hd };
assign dw_0[504] = dw_0_504[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_505 = { 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h3, 4'h5, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h3, 4'hc, 4'h0, 4'hf, 4'hc, 4'h1, 4'h0, 4'h1, 4'h5, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'hd, 4'h3, 4'h4, 4'hc };
assign dw_0[505] = dw_0_505[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_506 = { 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'hd, 4'hc, 4'h0, 4'hf, 4'h1, 4'hc, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'hf, 4'h0, 4'h4, 4'hd, 4'h4, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h7, 4'h3, 4'hd, 4'h3, 4'h3, 4'h0, 4'hd, 4'hc, 4'h1, 4'h5, 4'h3, 4'hc, 4'h0, 4'h5, 4'h0, 4'h3, 4'h3, 4'h3, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc };
assign dw_0[506] = dw_0_506[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_507 = { 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h7, 4'hc, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hf, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h1, 4'hd, 4'h4, 4'h3, 4'hd, 4'h0, 4'hf, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h5, 4'h7, 4'h0, 4'hf, 4'h0, 4'h0, 4'hd, 4'h3, 4'h4, 4'hd };
assign dw_0[507] = dw_0_507[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_508 = { 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h7, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'h1, 4'h4, 4'hd, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'hc, 4'h4, 4'h3, 4'h1, 4'h3, 4'hf, 4'h1, 4'h1, 4'h4, 4'h1, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h5, 4'h7, 4'h7, 4'hf, 4'h3, 4'h0, 4'hc, 4'h3, 4'h4, 4'hc };
assign dw_0[508] = dw_0_508[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_509 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'h7, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h1, 4'h0, 4'hd, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h0, 4'hd, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h3, 4'h1, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h5, 4'h7, 4'h3, 4'hf, 4'h0, 4'h0, 4'hd, 4'h3, 4'h4, 4'hc };
assign dw_0[509] = dw_0_509[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_510 = { 4'h1, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'h4, 4'hf, 4'h0, 4'hf, 4'h7, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h7, 4'hd, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'hf, 4'h3, 4'h1, 4'hd, 4'h0, 4'h1, 4'h0, 4'h3, 4'hd, 4'h3, 4'h5, 4'hc, 4'h7, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3, 4'h1, 4'h3, 4'h3, 4'hc, 4'h3, 4'h0, 4'hc, 4'h3, 4'h4, 4'hc };
assign dw_0[510] = dw_0_510[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_511 = { 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h7, 4'hd, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'hc, 4'h4, 4'hc, 4'h0, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'h0, 4'hd, 4'h4, 4'h0, 4'hd, 4'h0, 4'hf, 4'h5, 4'hd, 4'hc, 4'h1, 4'h4, 4'h3, 4'h1, 4'h3, 4'h5, 4'hc, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h5, 4'h3, 4'h4, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'hc };
assign dw_0[511] = dw_0_511[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_512 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'h3, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h0, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h5, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h1, 4'h0, 4'h0, 4'hd, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc };
assign dw_0[512] = dw_0_512[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_513 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hd, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'h3, 4'h3, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h5, 4'h0, 4'hd, 4'h5, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[513] = dw_0_513[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_514 = { 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'h4, 4'hc, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h7, 4'h5, 4'h3, 4'hc, 4'h1, 4'h0, 4'hf, 4'h3, 4'hf, 4'h1, 4'hc, 4'hc, 4'hd, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc };
assign dw_0[514] = dw_0_514[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_515 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h4, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h7, 4'h3, 4'h1, 4'h4, 4'hc, 4'hc, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h7, 4'h5, 4'hc, 4'hd, 4'h1, 4'h0, 4'hc, 4'h3, 4'hf, 4'h1, 4'hc, 4'hc, 4'h1, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'hf };
assign dw_0[515] = dw_0_515[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_516 = { 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hf, 4'hd, 4'h0, 4'h3, 4'hf, 4'h3, 4'h3, 4'h4, 4'h1, 4'hc, 4'hc, 4'h3, 4'h3, 4'h7, 4'h3, 4'h0, 4'h4, 4'hc, 4'hc, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'h7, 4'h5, 4'h7, 4'h1, 4'h1, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'hd, 4'hc, 4'h1, 4'h7, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf };
assign dw_0[516] = dw_0_516[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_517 = { 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h7, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h4, 4'h5, 4'h7, 4'hc, 4'hd, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc };
assign dw_0[517] = dw_0_517[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_518 = { 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'hd, 4'hc, 4'h3, 4'h3, 4'h7, 4'h3, 4'h0, 4'h4, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'hf, 4'h7, 4'h5, 4'h4, 4'h1, 4'h1, 4'h0, 4'h3, 4'h3, 4'hf, 4'hd, 4'h1, 4'hc, 4'h1, 4'h3, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h3, 4'hd, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc };
assign dw_0[518] = dw_0_518[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_519 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h1, 4'hc, 4'hc, 4'h3, 4'h3, 4'h7, 4'h3, 4'h0, 4'h4, 4'hd, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h3, 4'h5, 4'h3, 4'h0, 4'h5, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h3, 4'hc, 4'h0, 4'h7, 4'h3, 4'h3, 4'hf, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'hc, 4'hf };
assign dw_0[519] = dw_0_519[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_520 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h7, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h7, 4'h5, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc };
assign dw_0[520] = dw_0_520[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_521 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h5, 4'h3, 4'hc, 4'h5, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[521] = dw_0_521[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_522 = { 4'h3, 4'h3, 4'hc, 4'h3, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'hc, 4'h3, 4'h3, 4'h7, 4'h3, 4'h0, 4'h4, 4'hd, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h5, 4'h0, 4'h1, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'hd, 4'h0, 4'h0, 4'h7, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0 };
assign dw_0[522] = dw_0_522[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_523 = { 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'h7, 4'h3, 4'h1, 4'h4, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h4, 4'h3, 4'hc, 4'hd, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0 };
assign dw_0[523] = dw_0_523[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_524 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h4, 4'h1, 4'hc, 4'hc, 4'h0, 4'h3, 4'h7, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h4, 4'h3, 4'hd, 4'h1, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'h3, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc };
assign dw_0[524] = dw_0_524[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_525 = { 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h4, 4'h0, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'hf, 4'h4, 4'h5, 4'h7, 4'hc, 4'h5, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hd, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3 };
assign dw_0[525] = dw_0_525[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_526 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h7, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h5, 4'h3, 4'hc, 4'h5, 4'h0, 4'h0, 4'h3, 4'hf, 4'hd, 4'h0, 4'h0, 4'h1, 4'h3, 4'hf, 4'hc, 4'h0, 4'h7, 4'h0, 4'h3, 4'hc, 4'hc, 4'h5, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h4, 4'h3 };
assign dw_0[526] = dw_0_526[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_527 = { 4'h3, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h3, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h7, 4'h3, 4'h0, 4'h4, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h3, 4'h0, 4'h1, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h1, 4'h0, 4'hd, 4'h7, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'hd, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0 };
assign dw_0[527] = dw_0_527[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_528 = { 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'h4, 4'h3, 4'h3, 4'h1, 4'h3, 4'h5, 4'h3, 4'h5, 4'hd, 4'h1, 4'h1, 4'h5, 4'h3, 4'h3, 4'h5, 4'h4, 4'h1, 4'h4, 4'h0, 4'h4, 4'h4, 4'hd, 4'h0, 4'hd, 4'hf, 4'h7, 4'h3, 4'h5, 4'hc, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h5, 4'hd, 4'h1, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h7, 4'hd, 4'h0, 4'h7, 4'hc, 4'h4, 4'h0 };
assign dw_0[528] = dw_0_528[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_529 = { 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hd, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h5, 4'h3, 4'h4, 4'hc, 4'h1, 4'h5, 4'h1, 4'hf, 4'h4, 4'h4, 4'h0, 4'hd, 4'h1, 4'hc, 4'h0, 4'h0, 4'hd, 4'h0, 4'hd, 4'hf, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'hd, 4'h0, 4'hc, 4'h0, 4'h4, 4'hd, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1 };
assign dw_0[529] = dw_0_529[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_530 = { 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hd, 4'h7, 4'h3, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h5, 4'h7, 4'h4, 4'h0, 4'h1, 4'h5, 4'h1, 4'hf, 4'h0, 4'h4, 4'h4, 4'hd, 4'h5, 4'h0, 4'h0, 4'h7, 4'hd, 4'h0, 4'hd, 4'hf, 4'h3, 4'h0, 4'h4, 4'hc, 4'h1, 4'h1, 4'hc, 4'hc, 4'hc, 4'h1, 4'hd, 4'h1, 4'h0, 4'h5, 4'hc, 4'hc, 4'h0, 4'h1, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1 };
assign dw_0[530] = dw_0_530[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_531 = { 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'h7, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h7, 4'h5, 4'h3, 4'h4, 4'h3, 4'h1, 4'h1, 4'h0, 4'hf, 4'h4, 4'h5, 4'h4, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'hd, 4'h5, 4'hc, 4'hf, 4'h3, 4'h0, 4'h1, 4'hf, 4'hc, 4'h4, 4'hd, 4'h0, 4'h3, 4'h4, 4'hd, 4'hd, 4'h0, 4'h5, 4'hd, 4'hf, 4'hc, 4'h1, 4'hf, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0 };
assign dw_0[531] = dw_0_531[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_532 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'h7, 4'h7, 4'h3, 4'h3, 4'h0, 4'hc, 4'h4, 4'h5, 4'h3, 4'h4, 4'hf, 4'h1, 4'h1, 4'h0, 4'h3, 4'h4, 4'h4, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h7, 4'hd, 4'h5, 4'hc, 4'hf, 4'h0, 4'hf, 4'h1, 4'hf, 4'hd, 4'hd, 4'hc, 4'h0, 4'hd, 4'h0, 4'hd, 4'hc, 4'h0, 4'h4, 4'hc, 4'h3, 4'hc, 4'h1, 4'h3, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4 };
assign dw_0[532] = dw_0_532[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_533 = { 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5, 4'h3, 4'h4, 4'h3, 4'h1, 4'h1, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'hd, 4'h5, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'hc, 4'hf, 4'h3, 4'hc, 4'h1, 4'hf, 4'h1, 4'h0, 4'h1, 4'h0, 4'hc, 4'h5, 4'hd, 4'h1, 4'h0, 4'h4, 4'hc, 4'h0, 4'hc, 4'h5, 4'h3, 4'h0, 4'h3, 4'h1, 4'hf, 4'hf, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0 };
assign dw_0[533] = dw_0_533[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_534 = { 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'h4, 4'h5, 4'h3, 4'h5, 4'h3, 4'h1, 4'h5, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h4, 4'hc, 4'hf, 4'h3, 4'hf, 4'h1, 4'hf, 4'hc, 4'h0, 4'hc, 4'hc, 4'hc, 4'h4, 4'hd, 4'h1, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0 };
assign dw_0[534] = dw_0_534[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_535 = { 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'hd, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h7, 4'h5, 4'h3, 4'h4, 4'hf, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h7, 4'h4, 4'hd, 4'h0, 4'hc, 4'h0, 4'h3, 4'hd, 4'h1, 4'hc, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'hc, 4'hd, 4'h0, 4'hc, 4'hc, 4'h7, 4'hd, 4'h1, 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'hd, 4'h3, 4'hf, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0 };
assign dw_0[535] = dw_0_535[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_536 = { 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'h7, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h4, 4'h3, 4'h4, 4'hf, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'h4, 4'hd, 4'h0, 4'hc, 4'h0, 4'h3, 4'hd, 4'h1, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'hf, 4'hd, 4'hd, 4'h0, 4'h0, 4'h3, 4'h3, 4'hd, 4'h0, 4'h0, 4'h5, 4'hc, 4'h3, 4'h4, 4'h1, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'hf, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h4, 4'h1 };
assign dw_0[536] = dw_0_536[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_537 = { 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hd, 4'h4, 4'h4, 4'h3, 4'h3, 4'h3, 4'h5, 4'h7, 4'h4, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h4, 4'h4, 4'h4, 4'hd, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'hd, 4'hd, 4'h0, 4'h0, 4'h7, 4'hd, 4'h1, 4'h0, 4'h7, 4'hd, 4'h0, 4'h4, 4'h1, 4'h7, 4'h0, 4'h3, 4'h1, 4'hf, 4'hf, 4'h4, 4'h1, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0 };
assign dw_0[537] = dw_0_537[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_538 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'h7, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h3, 4'h4, 4'h0, 4'h1, 4'h4, 4'h1, 4'hf, 4'h4, 4'h4, 4'h4, 4'hd, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h3, 4'h4, 4'hd, 4'hc, 4'h7, 4'h1, 4'h3, 4'h0, 4'h3, 4'hd, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h4 };
assign dw_0[538] = dw_0_538[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_539 = { 4'h0, 4'hf, 4'hc, 4'h1, 4'h0, 4'h1, 4'h7, 4'h3, 4'hc, 4'hf, 4'h3, 4'h1, 4'h0, 4'h4, 4'h3, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'h7, 4'hc, 4'h1, 4'hc, 4'h3, 4'h3, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'h4, 4'hd, 4'hc, 4'h0, 4'h5, 4'hc, 4'hc, 4'h4, 4'h1, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4 };
assign dw_0[539] = dw_0_539[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_540 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h3, 4'h0, 4'h3, 4'h3, 4'h1, 4'h4, 4'h5, 4'h3, 4'h4, 4'hc, 4'h1, 4'h5, 4'h1, 4'h3, 4'h4, 4'h4, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'hd, 4'hc, 4'h0, 4'h5, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4 };
assign dw_0[540] = dw_0_540[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_541 = { 4'h3, 4'hc, 4'hc, 4'h1, 4'h0, 4'hc, 4'h7, 4'h4, 4'h4, 4'h0, 4'hf, 4'h4, 4'h4, 4'h4, 4'h3, 4'h5, 4'h0, 4'h1, 4'h5, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h7, 4'hd, 4'hd, 4'hc, 4'hf, 4'hf, 4'hc, 4'h4, 4'hc, 4'hd, 4'h1, 4'h0, 4'hc, 4'hc, 4'h4, 4'hd, 4'h0, 4'h0, 4'h5, 4'hd, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0 };
assign dw_0[541] = dw_0_541[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_542 = { 4'h3, 4'hd, 4'hc, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hf, 4'h0, 4'h5, 4'h1, 4'h3, 4'h4, 4'h4, 4'h0, 4'hc, 4'h1, 4'hc, 4'h0, 4'h7, 4'hd, 4'h1, 4'hd, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hd, 4'h1, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'h5, 4'hd, 4'h0, 4'h4, 4'h1, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0 };
assign dw_0[542] = dw_0_542[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_543 = { 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hd, 4'h7, 4'h4, 4'hf, 4'hf, 4'h3, 4'h1, 4'h0, 4'h5, 4'h3, 4'h4, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'h4, 4'h4, 4'h1, 4'h5, 4'hc, 4'h0, 4'h4, 4'hd, 4'h3, 4'hd, 4'hf, 4'h3, 4'h3, 4'h1, 4'h3, 4'h0, 4'hd, 4'h4, 4'hc, 4'h5, 4'h4, 4'hd, 4'hd, 4'h0, 4'h5, 4'hc, 4'hf, 4'h4, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'h5 };
assign dw_0[543] = dw_0_543[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_544 = { 4'h3, 4'h5, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'h0, 4'h1, 4'h5, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'hd, 4'h1, 4'h0, 4'h4, 4'h3, 4'h4, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'h1, 4'hc, 4'hd, 4'hd, 4'hf, 4'hc, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h5, 4'h3, 4'h0, 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'hc, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h5 };
assign dw_0[544] = dw_0_544[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_545 = { 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h5, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h7, 4'hc, 4'hc, 4'hc, 4'hd, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h4, 4'h4, 4'hd, 4'h0, 4'h1, 4'h0, 4'hd, 4'hd, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'hf, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h5 };
assign dw_0[545] = dw_0_545[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_546 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'h4, 4'hd, 4'h4, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h5, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'h4, 4'h5, 4'h0, 4'h5, 4'hc, 4'hd, 4'hd, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h7, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5 };
assign dw_0[546] = dw_0_546[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_547 = { 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h5, 4'h1, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h5, 4'h0, 4'h0, 4'h3, 4'h5, 4'hc, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'h1, 4'h3, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h3, 4'hd, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h5 };
assign dw_0[547] = dw_0_547[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_548 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h7, 4'h4, 4'h3, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'hd, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h5 };
assign dw_0[548] = dw_0_548[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_549 = { 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'hc, 4'h5, 4'h0, 4'hc, 4'h0, 4'h1, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'h4, 4'h5, 4'h1, 4'h0, 4'h4, 4'h0, 4'hd, 4'h1, 4'h3, 4'hc, 4'hf, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5 };
assign dw_0[549] = dw_0_549[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_550 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'hd, 4'h5, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hd, 4'h5, 4'h4, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'hc, 4'hd, 4'hd, 4'h3, 4'hc, 4'hf, 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5 };
assign dw_0[550] = dw_0_550[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_551 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h7, 4'hc, 4'h5, 4'h0, 4'h1, 4'h5, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'h1, 4'h4, 4'h0, 4'h7, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'h1, 4'h0, 4'hc, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'hc, 4'h4, 4'h0, 4'h0, 4'h7, 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5 };
assign dw_0[551] = dw_0_551[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_552 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h1, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h5 };
assign dw_0[552] = dw_0_552[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_553 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'h3, 4'h1, 4'h0, 4'hd, 4'h4, 4'h0, 4'h5, 4'h0, 4'h1, 4'h7, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc, 4'h1, 4'h5, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h5, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'hd, 4'h1, 4'h3, 4'h0, 4'hc, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'hd, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h5 };
assign dw_0[553] = dw_0_553[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_554 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'h1, 4'h4, 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'hd, 4'hd, 4'h3, 4'h0, 4'hf, 4'h3, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hd, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5 };
assign dw_0[554] = dw_0_554[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_555 = { 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'h0, 4'h0, 4'hf, 4'hc, 4'hd, 4'h4, 4'h4, 4'h0, 4'h7, 4'h4, 4'h4, 4'h0, 4'hd, 4'h1, 4'h0, 4'h4, 4'h0, 4'hd, 4'hd, 4'hf, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5 };
assign dw_0[555] = dw_0_555[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_556 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h7, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h4, 4'hd, 4'h5, 4'h0, 4'h1, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'h5, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'h5, 4'h1, 4'h0, 4'h4, 4'hc, 4'hd, 4'hd, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5 };
assign dw_0[556] = dw_0_556[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_557 = { 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h1, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'hc, 4'h4, 4'h1, 4'h1, 4'h3, 4'h4, 4'h0, 4'hd, 4'hd, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h7, 4'h1, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h5 };
assign dw_0[557] = dw_0_557[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_558 = { 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hd, 4'hc, 4'h7, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hd, 4'h5, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'hd, 4'hd, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h7, 4'h1, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h5 };
assign dw_0[558] = dw_0_558[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_559 = { 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h3, 4'h0, 4'hc, 4'hf, 4'hc, 4'hd, 4'h5, 4'h4, 4'h0, 4'h3, 4'h4, 4'hc, 4'h4, 4'h4, 4'hd, 4'h0, 4'h5, 4'h0, 4'hd, 4'hd, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h7, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'hf, 4'h0, 4'h4, 4'h5 };
assign dw_0[559] = dw_0_559[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_560 = { 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h1, 4'h3, 4'h4, 4'hc, 4'h0, 4'h1, 4'h3, 4'hf, 4'h3, 4'hc, 4'h1, 4'h0, 4'h3, 4'hd, 4'h0, 4'h3, 4'hc, 4'hf, 4'h4, 4'h0, 4'hd, 4'h4, 4'h0, 4'hd, 4'hd, 4'hd, 4'h7, 4'h4, 4'hf, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc, 4'h7, 4'hc, 4'hf, 4'hd, 4'h4, 4'h0, 4'h0, 4'h7, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h4 };
assign dw_0[560] = dw_0_560[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_561 = { 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h7, 4'h4, 4'h0, 4'h0, 4'hf, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'h7, 4'h5, 4'hf, 4'h0, 4'h4, 4'h0, 4'hd, 4'h3, 4'hf, 4'hc, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'hf, 4'hc, 4'h4, 4'h0, 4'h0, 4'h7, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h4 };
assign dw_0[561] = dw_0_561[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_562 = { 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h1, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h7, 4'h0, 4'hf, 4'h0, 4'h1, 4'hc, 4'h5, 4'h0, 4'hf, 4'hc, 4'hf, 4'hd, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'hd, 4'hc, 4'h4, 4'h0, 4'h0, 4'h7, 4'h4, 4'h5, 4'h3, 4'h5, 4'h0, 4'h7, 4'h3, 4'h0, 4'h7 };
assign dw_0[562] = dw_0_562[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_563 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'hd, 4'h3, 4'h4, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc, 4'h3, 4'hc, 4'hf, 4'hd, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'hf, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3 };
assign dw_0[563] = dw_0_563[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_564 = { 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'hf, 4'h1, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'h3, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'h3, 4'h4, 4'hc, 4'h3, 4'hc, 4'hf, 4'hd, 4'h3, 4'hf, 4'h0, 4'h7, 4'h3, 4'h0, 4'hd, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[564] = dw_0_564[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_565 = { 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h5, 4'h4, 4'h3, 4'h1, 4'hf, 4'h4, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'h5, 4'h0, 4'hc, 4'h3, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'hd, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'hc, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3 };
assign dw_0[565] = dw_0_565[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_566 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h3, 4'h4, 4'h7, 4'h0, 4'h1, 4'h3, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h7, 4'h1, 4'hf, 4'h0, 4'h1, 4'h3, 4'h1, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'h4, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'hd, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[566] = dw_0_566[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_567 = { 4'h1, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'hd, 4'hc, 4'h3, 4'h4, 4'hf, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'h7, 4'h4, 4'h7, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[567] = dw_0_567[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_568 = { 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h1, 4'hf, 4'h5, 4'h4, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h3, 4'hc, 4'h3, 4'h4, 4'h3, 4'h0, 4'h4, 4'h4, 4'hf, 4'h1, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'hd, 4'hc, 4'h0, 4'h7, 4'h3, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0 };
assign dw_0[568] = dw_0_568[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_569 = { 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'hc, 4'hc, 4'h1, 4'h0, 4'hd, 4'h1, 4'h3, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'hc, 4'h7, 4'h4, 4'hf, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'h5, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0 };
assign dw_0[569] = dw_0_569[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_570 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h4, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'h3, 4'hd, 4'hc, 4'h0, 4'h3, 4'hd, 4'h5, 4'h7, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h7, 4'h4, 4'hc, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc, 4'h3, 4'hc, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'hc, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4 };
assign dw_0[570] = dw_0_570[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_571 = { 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h7, 4'h5, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'hc, 4'hf, 4'hc, 4'h4, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[571] = dw_0_571[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_572 = { 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h7, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h1, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'hc, 4'h7, 4'h4, 4'hf, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'h1, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3 };
assign dw_0[572] = dw_0_572[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_573 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hd, 4'h0, 4'hc, 4'h0, 4'h7, 4'h3, 4'h3, 4'h4, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3 };
assign dw_0[573] = dw_0_573[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_574 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'hc, 4'hf, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'h4, 4'hc, 4'hc, 4'h4, 4'hc, 4'hc, 4'h5, 4'hc, 4'h7, 4'h4, 4'hf, 4'h0, 4'h5, 4'hd, 4'h0, 4'h3, 4'h3, 4'hc, 4'hf, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'hd, 4'h0, 4'h7, 4'h4, 4'h0, 4'h3 };
assign dw_0[574] = dw_0_574[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_575 = { 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h5, 4'h4, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'hd, 4'h1, 4'h0, 4'hc, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h4, 4'hf, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'h1, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'h5, 4'h5, 4'h1, 4'h1, 4'h0, 4'h7, 4'h0, 4'hc, 4'h0 };
assign dw_0[575] = dw_0_575[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_576 = { 4'hc, 4'h7, 4'h0, 4'h1, 4'h0, 4'h4, 4'h5, 4'h7, 4'h4, 4'h1, 4'hc, 4'h4, 4'h3, 4'h4, 4'h4, 4'h3, 4'hc, 4'h1, 4'hc, 4'h5, 4'hc, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'h3, 4'hd, 4'h4, 4'h4, 4'hc, 4'h7, 4'hd, 4'h4, 4'hc, 4'h3, 4'h1, 4'h5, 4'h0, 4'hc, 4'h5, 4'h5, 4'hf, 4'h1, 4'h3, 4'h0, 4'h4, 4'hf, 4'h0, 4'h0, 4'hd, 4'hf, 4'h0, 4'hf, 4'h5, 4'h4, 4'h3 };
assign dw_0[576] = dw_0_576[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_577 = { 4'h1, 4'h7, 4'hc, 4'h1, 4'h0, 4'h7, 4'h7, 4'h7, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'h1, 4'hf, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'hc, 4'hc, 4'h3, 4'hc, 4'hd, 4'h3, 4'h7, 4'h3, 4'h1, 4'h5, 4'h0, 4'h0, 4'h7, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'h1, 4'hd, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'hd, 4'h3, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0 };
assign dw_0[577] = dw_0_577[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_578 = { 4'h1, 4'h7, 4'hc, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'hc, 4'h1, 4'hc, 4'h7, 4'h0, 4'h7, 4'h4, 4'h0, 4'hf, 4'h0, 4'hc, 4'hd, 4'hd, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'h7, 4'h0, 4'h4, 4'h4, 4'h7, 4'h7, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'h1, 4'h1, 4'h4, 4'hf, 4'h0, 4'hf, 4'h0, 4'h3, 4'hf, 4'h0, 4'h3, 4'hd, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0 };
assign dw_0[578] = dw_0_578[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_579 = { 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'hc, 4'h0, 4'h1, 4'h7, 4'h7, 4'h3, 4'h4, 4'h0, 4'hf, 4'h0, 4'hc, 4'h1, 4'hc, 4'h0, 4'hf, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'hc, 4'h3, 4'h7, 4'h3, 4'h3, 4'h5, 4'h4, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'h1, 4'h1, 4'hd, 4'h0, 4'h4, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0 };
assign dw_0[579] = dw_0_579[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_580 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'h7, 4'h3, 4'h4, 4'h4, 4'hf, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h7, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'h3, 4'h4, 4'h4, 4'h1, 4'hc, 4'h0, 4'h1, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h4, 4'hc, 4'h0 };
assign dw_0[580] = dw_0_580[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_581 = { 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'hd, 4'h0, 4'h3, 4'h7, 4'h4, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'hd, 4'h4, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h3, 4'h7, 4'h3, 4'h0, 4'h7, 4'h4, 4'h0, 4'h7, 4'h5, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'hf, 4'h0, 4'hf, 4'h0, 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h0 };
assign dw_0[581] = dw_0_581[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_582 = { 4'h1, 4'h7, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h7, 4'h4, 4'hf, 4'h0, 4'hc, 4'h3, 4'hc, 4'h7, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h3, 4'h3, 4'h4, 4'h3, 4'h0, 4'h7, 4'h5, 4'h4, 4'h0, 4'h4, 4'h4, 4'hc, 4'h1, 4'h1, 4'h0, 4'h4, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0 };
assign dw_0[582] = dw_0_582[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_583 = { 4'h0, 4'h7, 4'hc, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h7, 4'h0, 4'hf, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h7, 4'h5, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h5, 4'h0, 4'h0 };
assign dw_0[583] = dw_0_583[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_584 = { 4'h0, 4'h7, 4'hc, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'hf, 4'h1, 4'hd, 4'h7, 4'h3, 4'h3, 4'h4, 4'h4, 4'h3, 4'h3, 4'h1, 4'h3, 4'h3, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h7, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'h7, 4'h5, 4'h0, 4'h0, 4'h7, 4'h7, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc, 4'h4, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc };
assign dw_0[584] = dw_0_584[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_585 = { 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h3, 4'hc, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h7, 4'h4, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'h4, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'hc, 4'hc, 4'h3, 4'h3, 4'h3, 4'h5, 4'h0, 4'h0, 4'h7, 4'h1, 4'h4, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h5, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0 };
assign dw_0[585] = dw_0_585[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_586 = { 4'h1, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h1, 4'h1, 4'h3, 4'hd, 4'h0, 4'hc, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h7, 4'h4, 4'h4, 4'h1, 4'h3, 4'h3, 4'h1, 4'h0, 4'hc, 4'h0, 4'h1, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0 };
assign dw_0[586] = dw_0_586[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_587 = { 4'hd, 4'h7, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h7, 4'h3, 4'h4, 4'h3, 4'h4, 4'h4, 4'h7, 4'h7, 4'h5, 4'h4, 4'h1, 4'h7, 4'h3, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'hf, 4'h1, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0 };
assign dw_0[587] = dw_0_587[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_588 = { 4'hd, 4'h7, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h4, 4'h5, 4'h0, 4'hc, 4'hc, 4'h7, 4'hc, 4'hc, 4'h0, 4'h3, 4'h7, 4'h0, 4'h1, 4'h4, 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h4, 4'hf, 4'h1, 4'hf, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h5, 4'h0, 4'h0 };
assign dw_0[588] = dw_0_588[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_589 = { 4'hc, 4'h7, 4'h0, 4'h1, 4'h0, 4'h7, 4'h4, 4'h3, 4'hc, 4'h1, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h1, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3 };
assign dw_0[589] = dw_0_589[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_590 = { 4'hd, 4'h7, 4'h0, 4'h1, 4'h0, 4'h7, 4'h4, 4'hf, 4'hc, 4'hd, 4'hf, 4'h7, 4'h0, 4'h3, 4'h4, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h7, 4'h3, 4'h3, 4'h5, 4'h7, 4'h3, 4'h7, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h5, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'hd, 4'h0, 4'hf, 4'h4, 4'h0, 4'h3 };
assign dw_0[590] = dw_0_590[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_591 = { 4'h1, 4'h7, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'hf, 4'hf, 4'h1, 4'hc, 4'h7, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h7, 4'h3, 4'hd, 4'hc, 4'h7, 4'h7, 4'h1, 4'h4, 4'h4, 4'h0, 4'h7, 4'hd, 4'h0, 4'hd, 4'h3, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h1, 4'hc, 4'h1, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hd, 4'h3, 4'h0, 4'h3, 4'h5, 4'hc, 4'h3 };
assign dw_0[591] = dw_0_591[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_592 = { 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h7, 4'hd, 4'h0, 4'h7, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h1, 4'hc, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'h4, 4'hc, 4'hd, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h3 };
assign dw_0[592] = dw_0_592[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_593 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'hf, 4'h3, 4'hd, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h4, 4'h0, 4'hd, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h3, 4'h7, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3 };
assign dw_0[593] = dw_0_593[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_594 = { 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h4, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'hc, 4'hd, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3 };
assign dw_0[594] = dw_0_594[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_595 = { 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h3, 4'hd, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h3, 4'h7, 4'hd, 4'h0, 4'h4, 4'hc, 4'h1, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hc, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3 };
assign dw_0[595] = dw_0_595[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_596 = { 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h3, 4'h0, 4'hd, 4'h0, 4'h7, 4'h0, 4'h1, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h4, 4'h0, 4'h3, 4'h4, 4'hd, 4'h0, 4'h0, 4'hc, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'hc, 4'h3 };
assign dw_0[596] = dw_0_596[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_597 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'hc, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h3, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3 };
assign dw_0[597] = dw_0_597[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_598 = { 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'h4, 4'h3, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0 };
assign dw_0[598] = dw_0_598[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_599 = { 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'hd, 4'h0, 4'hf, 4'h3, 4'h1, 4'h0, 4'h4, 4'h3, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h7, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3 };
assign dw_0[599] = dw_0_599[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_600 = { 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h7, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0 };
assign dw_0[600] = dw_0_600[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_601 = { 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h3, 4'hd, 4'hf, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'h0, 4'hf, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'hf, 4'h1, 4'h0, 4'h4, 4'h7, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'hd, 4'h3, 4'h0, 4'h3 };
assign dw_0[601] = dw_0_601[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_602 = { 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3 };
assign dw_0[602] = dw_0_602[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_603 = { 4'hc, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h5, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3 };
assign dw_0[603] = dw_0_603[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_604 = { 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h4, 4'hd, 4'h3, 4'h3, 4'h4, 4'hd, 4'h3, 4'h7, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hd, 4'h4, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0 };
assign dw_0[604] = dw_0_604[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_605 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'hd, 4'h3, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'hf, 4'hd, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'hf, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3 };
assign dw_0[605] = dw_0_605[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_606 = { 4'h1, 4'h5, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'hf, 4'h0, 4'hd, 4'h0, 4'h4, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h4, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'hf, 4'hd, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'hf, 4'h0, 4'hd, 4'h0, 4'hc, 4'h3 };
assign dw_0[606] = dw_0_606[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_607 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h1, 4'hf, 4'h0, 4'hd, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'hc, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h4, 4'h4, 4'h1, 4'hd, 4'h0, 4'h4, 4'hc, 4'hc, 4'h4, 4'h0, 4'h3, 4'h1, 4'h1, 4'h3, 4'h5, 4'hc, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3 };
assign dw_0[607] = dw_0_607[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_608 = { 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h4, 4'h3, 4'h3, 4'h4, 4'h0, 4'h4, 4'hd, 4'h3, 4'hc, 4'hf, 4'h3, 4'h1, 4'h1, 4'hc, 4'h3, 4'h1, 4'h0, 4'h4, 4'h5, 4'h4, 4'hc, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h7, 4'hc, 4'h5, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc };
assign dw_0[608] = dw_0_608[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_609 = { 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'hf, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'hd, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'hd, 4'hc, 4'h7, 4'hc, 4'h4, 4'h0, 4'h3, 4'h5, 4'hc, 4'h0, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hd };
assign dw_0[609] = dw_0_609[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_610 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h4, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'hd, 4'hc, 4'h7, 4'h0, 4'h1, 4'hc, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'hc };
assign dw_0[610] = dw_0_610[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_611 = { 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hd, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h4, 4'hd, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'hc, 4'hf, 4'h3, 4'h0, 4'h1, 4'hc, 4'h3, 4'h5, 4'h0, 4'h4, 4'h4, 4'h7, 4'hc, 4'h0, 4'h0, 4'h5, 4'hc, 4'hc, 4'hf, 4'h7, 4'h1, 4'h0, 4'h3, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'hc };
assign dw_0[611] = dw_0_611[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_612 = { 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h3, 4'h4, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h1, 4'hc, 4'h3, 4'hc, 4'hc, 4'h4, 4'h3, 4'h1, 4'hc, 4'h3, 4'h5, 4'h0, 4'h4, 4'h5, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h7, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'hc };
assign dw_0[612] = dw_0_612[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_613 = { 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'hc, 4'h7, 4'h3, 4'h0, 4'hc, 4'h3, 4'hd, 4'h4, 4'h4, 4'h4, 4'h0, 4'hf, 4'h1, 4'h3, 4'h4, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3, 4'hf, 4'h1, 4'h0, 4'hc, 4'h3, 4'h4, 4'hc };
assign dw_0[613] = dw_0_613[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_614 = { 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h3, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'hc, 4'h3, 4'h3, 4'h1, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h3, 4'h0, 4'h0, 4'h5, 4'hf, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hc };
assign dw_0[614] = dw_0_614[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_615 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h4, 4'h4, 4'hc, 4'h0, 4'h7, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'hc, 4'h7, 4'h3, 4'h1, 4'hc, 4'h3, 4'hd, 4'h4, 4'h4, 4'h4, 4'h4, 4'hc, 4'h1, 4'h0, 4'h1, 4'hc, 4'h1, 4'h3, 4'h3, 4'h1, 4'h0, 4'h3, 4'h5, 4'h0, 4'h3, 4'hf, 4'h1, 4'h0, 4'h0, 4'hf, 4'h4, 4'hc };
assign dw_0[615] = dw_0_615[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_616 = { 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'hd, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h7, 4'h0, 4'h1, 4'hc, 4'h3, 4'h1, 4'h1, 4'h4, 4'h4, 4'h7, 4'hf, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h1, 4'hc, 4'h4, 4'hc };
assign dw_0[616] = dw_0_616[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_617 = { 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h3, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'hd, 4'h3, 4'hc, 4'hc, 4'h7, 4'h0, 4'hd, 4'hc, 4'hf, 4'h1, 4'h4, 4'h4, 4'h4, 4'h4, 4'h3, 4'h1, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc, 4'h7, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd };
assign dw_0[617] = dw_0_617[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_618 = { 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'hd, 4'h4, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'hf, 4'h7, 4'h0, 4'h1, 4'hc, 4'h3, 4'h1, 4'h5, 4'h0, 4'h4, 4'h4, 4'h3, 4'h1, 4'h0, 4'h5, 4'hd, 4'h0, 4'h7, 4'h3, 4'h1, 4'h0, 4'h3, 4'h5, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc };
assign dw_0[618] = dw_0_618[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_619 = { 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'h4, 4'hd, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc, 4'hf, 4'h7, 4'h0, 4'h1, 4'h0, 4'h7, 4'h5, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'hc, 4'h3, 4'h0, 4'hc, 4'h3, 4'h4, 4'hc };
assign dw_0[619] = dw_0_619[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_620 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'hd, 4'h4, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'h1, 4'h1, 4'h4, 4'h5, 4'h4, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h7, 4'h1, 4'h0, 4'h3, 4'h5, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc };
assign dw_0[620] = dw_0_620[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_621 = { 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'h5, 4'hc, 4'h7, 4'hd, 4'hf, 4'h7, 4'h0, 4'h1, 4'hc, 4'h3, 4'h5, 4'h1, 4'h0, 4'h5, 4'h7, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc };
assign dw_0[621] = dw_0_621[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_622 = { 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hc, 4'h1, 4'h0, 4'hf, 4'h0, 4'h3, 4'h1, 4'hf, 4'h4, 4'h1, 4'h0, 4'h1, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h3, 4'hc, 4'hc, 4'h7, 4'h1, 4'h5, 4'hc, 4'h7, 4'h5, 4'h1, 4'h0, 4'h5, 4'h0, 4'hc, 4'h1, 4'h3, 4'h1, 4'h0, 4'hc, 4'h3, 4'h3, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'hc };
assign dw_0[622] = dw_0_622[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_623 = { 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hd, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'h3, 4'hd, 4'h3, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'hf, 4'h0, 4'h0, 4'h5, 4'hd, 4'h3, 4'hd, 4'hc, 4'h7, 4'h1, 4'h1, 4'h0, 4'h7, 4'h5, 4'hc, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h5, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hc };
assign dw_0[623] = dw_0_623[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_624 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h3, 4'hc, 4'hc, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'h3, 4'h3, 4'hf, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'hf, 4'h1, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'hd, 4'hc, 4'h4, 4'h4, 4'h3, 4'h0, 4'hd, 4'h0, 4'h1, 4'hc, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h3, 4'hc, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'hf, 4'h4, 4'h0 };
assign dw_0[624] = dw_0_624[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_625 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h3, 4'hd, 4'hc, 4'h4, 4'h0, 4'h0, 4'h5, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hf };
assign dw_0[625] = dw_0_625[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_626 = { 4'hc, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'hf, 4'hc, 4'h4, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h7, 4'h3, 4'h0, 4'h0, 4'h7, 4'h0, 4'hf, 4'h1, 4'h0, 4'hc, 4'h0, 4'hd, 4'h5, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hf, 4'h4, 4'h0 };
assign dw_0[626] = dw_0_626[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_627 = { 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h1, 4'h3, 4'h0, 4'hd, 4'h0, 4'h3, 4'hc, 4'h1, 4'h4, 4'h0, 4'h3, 4'h4, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h7, 4'h5, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0 };
assign dw_0[627] = dw_0_627[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_628 = { 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h7, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'hc, 4'h4, 4'h4, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0 };
assign dw_0[628] = dw_0_628[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_629 = { 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'hf, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'h4, 4'h4, 4'hc, 4'h5, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h7, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0 };
assign dw_0[629] = dw_0_629[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_630 = { 4'hc, 4'h1, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3, 4'hc, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h0, 4'hd, 4'h1, 4'h4, 4'h0, 4'h3, 4'h4, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc };
assign dw_0[630] = dw_0_630[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_631 = { 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h4, 4'h3, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hd, 4'h4, 4'h4, 4'hc, 4'h0, 4'h4, 4'h3, 4'h3, 4'h4, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h7, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[631] = dw_0_631[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_632 = { 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'hf, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[632] = dw_0_632[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_633 = { 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'h4, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[633] = dw_0_633[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_634 = { 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'hc, 4'h4, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[634] = dw_0_634[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_635 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hd, 4'h0, 4'hc, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0 };
assign dw_0[635] = dw_0_635[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_636 = { 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hc, 4'hc, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hd, 4'h1, 4'h4, 4'h4, 4'hf, 4'h4, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3 };
assign dw_0[636] = dw_0_636[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_637 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h4, 4'h3, 4'hf, 4'hc, 4'hd, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h1, 4'hd, 4'h0, 4'hc, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h5, 4'hc, 4'h0, 4'h4, 4'hf, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h4, 4'h0 };
assign dw_0[637] = dw_0_637[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_638 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h3, 4'hc, 4'hc, 4'h4, 4'h0, 4'h3, 4'h5, 4'hd, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h7, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0 };
assign dw_0[638] = dw_0_638[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_639 = { 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h4, 4'hc, 4'h0, 4'h4, 4'h4, 4'h3, 4'h5, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h4, 4'h4, 4'h1, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hf, 4'h0, 4'h0 };
assign dw_0[639] = dw_0_639[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_640 = { 4'h3, 4'h1, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'hf, 4'h3, 4'hd, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h3, 4'h3, 4'h7, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h3, 4'h5, 4'hf, 4'h4, 4'hd, 4'hc, 4'h4, 4'h1, 4'h7, 4'h0, 4'hc, 4'h0, 4'h5, 4'hc, 4'h3, 4'hf, 4'h3, 4'h7, 4'h0, 4'h0, 4'hd, 4'hf, 4'hd, 4'h3, 4'h3, 4'h0, 4'hf, 4'hf, 4'h4, 4'h0 };
assign dw_0[640] = dw_0_640[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_641 = { 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h1, 4'h5, 4'h3, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h4, 4'hf, 4'h4, 4'h5, 4'hf, 4'h0, 4'h5, 4'hc, 4'h0, 4'hd, 4'hf, 4'h4, 4'h0, 4'h4, 4'h1, 4'hd, 4'h0, 4'h5, 4'hc, 4'hf, 4'h3, 4'h3, 4'h7, 4'h0, 4'h3, 4'h1, 4'hc, 4'hd, 4'hf, 4'h3, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0 };
assign dw_0[641] = dw_0_641[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_642 = { 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'hd, 4'h4, 4'h5, 4'h3, 4'hf, 4'h3, 4'hd, 4'h4, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h3, 4'h3, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h5, 4'hf, 4'h0, 4'h1, 4'hf, 4'hc, 4'hd, 4'h3, 4'h4, 4'h0, 4'h4, 4'hd, 4'hd, 4'h0, 4'h5, 4'hc, 4'hf, 4'hf, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'hc, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0 };
assign dw_0[642] = dw_0_642[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_643 = { 4'hf, 4'h1, 4'hc, 4'h3, 4'h0, 4'hc, 4'h4, 4'h5, 4'h3, 4'hf, 4'h0, 4'hc, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h3, 4'h3, 4'h0, 4'hd, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'hc, 4'h1, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h1, 4'hf, 4'hc, 4'hd, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'h4, 4'hc, 4'h3, 4'hf, 4'hc, 4'h7, 4'h0, 4'h3, 4'hd, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3 };
assign dw_0[643] = dw_0_643[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_644 = { 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h3, 4'hf, 4'h1, 4'h0, 4'h4, 4'h5, 4'hc, 4'h7, 4'h0, 4'h0, 4'h5, 4'h3, 4'h3, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h3, 4'h4, 4'h4, 4'hc, 4'h3, 4'h1, 4'hf, 4'hc, 4'hd, 4'h0, 4'h4, 4'h0, 4'h7, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h7, 4'h0, 4'hf, 4'hd, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h3 };
assign dw_0[644] = dw_0_644[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_645 = { 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hd, 4'h4, 4'h5, 4'hf, 4'hf, 4'h0, 4'hd, 4'h4, 4'h1, 4'hd, 4'h0, 4'h3, 4'h3, 4'h5, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h7, 4'h1, 4'hf, 4'h0, 4'h1, 4'hf, 4'h0, 4'hd, 4'h3, 4'h4, 4'h0, 4'h7, 4'hf, 4'hd, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'h3, 4'h7, 4'h0, 4'hf, 4'h1, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0 };
assign dw_0[645] = dw_0_645[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_646 = { 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h4, 4'h5, 4'hf, 4'hf, 4'h3, 4'hd, 4'h4, 4'h1, 4'hd, 4'h0, 4'h3, 4'h3, 4'h5, 4'h3, 4'h3, 4'h4, 4'h1, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h7, 4'h4, 4'hf, 4'h0, 4'h1, 4'hf, 4'hc, 4'hd, 4'h0, 4'h4, 4'h4, 4'h7, 4'hc, 4'hd, 4'h0, 4'h5, 4'h0, 4'h3, 4'hf, 4'h3, 4'h7, 4'h0, 4'h3, 4'h1, 4'hc, 4'hd, 4'hc, 4'h0, 4'h0, 4'h1, 4'hf, 4'h4, 4'h0 };
assign dw_0[646] = dw_0_646[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_647 = { 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h5, 4'h3, 4'hf, 4'h3, 4'hd, 4'h4, 4'h5, 4'hc, 4'h0, 4'h3, 4'h3, 4'h5, 4'h3, 4'h3, 4'h0, 4'hd, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'hf, 4'hc, 4'hf, 4'h7, 4'h0, 4'hf, 4'h0, 4'h1, 4'hf, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h0, 4'h4, 4'hc, 4'h3, 4'hf, 4'hc, 4'h7, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'h0 };
assign dw_0[647] = dw_0_647[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_648 = { 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h5, 4'h4, 4'h3, 4'hf, 4'h0, 4'hd, 4'h4, 4'h5, 4'hf, 4'h3, 4'h3, 4'h0, 4'h5, 4'h3, 4'h3, 4'h4, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h3, 4'h7, 4'h4, 4'hf, 4'h3, 4'h1, 4'hf, 4'h1, 4'hd, 4'hc, 4'h4, 4'hc, 4'h7, 4'h0, 4'hc, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'hc, 4'h7, 4'hc, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0 };
assign dw_0[648] = dw_0_648[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_649 = { 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'h5, 4'h3, 4'hf, 4'h3, 4'hc, 4'h4, 4'h5, 4'hd, 4'h3, 4'h0, 4'h3, 4'h5, 4'h3, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h5, 4'hc, 4'h3, 4'h4, 4'hf, 4'h0, 4'h1, 4'hf, 4'h1, 4'hd, 4'h1, 4'h4, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h5, 4'hc, 4'h3, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0 };
assign dw_0[649] = dw_0_649[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_650 = { 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h5, 4'h3, 4'hf, 4'h3, 4'hd, 4'h4, 4'h1, 4'hd, 4'h0, 4'h4, 4'h3, 4'h4, 4'h3, 4'h3, 4'h0, 4'hd, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'h1, 4'hf, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h5, 4'hc, 4'h3, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h4, 4'h3 };
assign dw_0[650] = dw_0_650[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_651 = { 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hd, 4'h4, 4'h5, 4'h3, 4'hf, 4'h3, 4'hd, 4'h4, 4'h1, 4'hd, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h3, 4'h4, 4'hd, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'h7, 4'h4, 4'hf, 4'h0, 4'h1, 4'hf, 4'hc, 4'hd, 4'h0, 4'h4, 4'h1, 4'h7, 4'h0, 4'hd, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h3, 4'h7, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'h4 };
assign dw_0[651] = dw_0_651[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_652 = { 4'h3, 4'hd, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h5, 4'h3, 4'hf, 4'hf, 4'hd, 4'h4, 4'h1, 4'hc, 4'h4, 4'h3, 4'h0, 4'h5, 4'h3, 4'h7, 4'h4, 4'hd, 4'hc, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'hf, 4'h4, 4'h5, 4'hf, 4'h0, 4'h1, 4'hf, 4'hc, 4'hd, 4'h0, 4'h4, 4'h1, 4'h7, 4'h0, 4'hc, 4'h0, 4'h5, 4'h1, 4'hf, 4'h3, 4'h3, 4'h7, 4'h0, 4'h3, 4'h1, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h4, 4'hf };
assign dw_0[652] = dw_0_652[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_653 = { 4'h3, 4'h1, 4'hc, 4'h0, 4'h0, 4'hd, 4'h0, 4'h5, 4'h0, 4'hf, 4'h3, 4'hd, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h3, 4'h3, 4'h4, 4'h1, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h4, 4'h5, 4'hf, 4'h3, 4'h1, 4'hf, 4'hc, 4'hd, 4'hc, 4'h0, 4'h0, 4'h7, 4'hc, 4'hd, 4'h0, 4'h5, 4'hc, 4'h3, 4'h3, 4'hc, 4'h7, 4'h0, 4'h0, 4'hd, 4'hf, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0 };
assign dw_0[653] = dw_0_653[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_654 = { 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h3, 4'h3, 4'h4, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'h4, 4'h4, 4'hf, 4'h0, 4'h1, 4'hf, 4'hc, 4'hd, 4'hf, 4'h4, 4'h0, 4'h7, 4'hc, 4'hc, 4'h0, 4'h4, 4'hc, 4'h3, 4'h3, 4'hf, 4'h7, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h4, 4'h0 };
assign dw_0[654] = dw_0_654[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_655 = { 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hc, 4'h4, 4'h5, 4'hf, 4'hf, 4'h3, 4'hd, 4'h0, 4'h5, 4'h0, 4'h5, 4'h0, 4'h0, 4'h5, 4'h3, 4'h3, 4'h0, 4'h1, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'hf, 4'h4, 4'h1, 4'h0, 4'h3, 4'h1, 4'hf, 4'hd, 4'hd, 4'h3, 4'h0, 4'h5, 4'h4, 4'hc, 4'hd, 4'h0, 4'h5, 4'hc, 4'hf, 4'h3, 4'h0, 4'h7, 4'h0, 4'h3, 4'h1, 4'h3, 4'h4, 4'h3, 4'h3, 4'h0, 4'hc, 4'hf, 4'h4, 4'h5 };
assign dw_0[655] = dw_0_655[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_656 = { 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h4, 4'hd, 4'hf, 4'h0, 4'hf, 4'h0, 4'hd, 4'hd, 4'h0, 4'h1, 4'h3, 4'h3, 4'hd, 4'h3, 4'hc, 4'h1, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h5, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'h1, 4'hc, 4'h0, 4'h7, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h1, 4'hf, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'h0, 4'hd, 4'h7, 4'h0, 4'hd, 4'h0, 4'h0, 4'hf };
assign dw_0[656] = dw_0_656[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_657 = { 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h1, 4'hc, 4'hd, 4'h0, 4'h1, 4'hd, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'hf, 4'hc, 4'h4, 4'hc, 4'h4, 4'h1, 4'h4, 4'h0, 4'hc, 4'h3, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'hc, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h1, 4'hd, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h7, 4'h0, 4'hc };
assign dw_0[657] = dw_0_657[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_658 = { 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'hc, 4'hd, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'h7, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h1, 4'h7, 4'h0, 4'hc, 4'h3, 4'h1, 4'h0, 4'h4, 4'h3, 4'h4, 4'hc, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0 };
assign dw_0[658] = dw_0_658[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_659 = { 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'hd, 4'hf, 4'h4, 4'h3, 4'h7, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'hd, 4'h4, 4'h0, 4'h5, 4'h7, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h5, 4'h1, 4'h7, 4'hc, 4'hc, 4'h3, 4'h5, 4'hc, 4'h4, 4'h7, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[659] = dw_0_659[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_660 = { 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h7, 4'h3, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'hd, 4'h0, 4'h1, 4'hc, 4'h7, 4'h0, 4'h3, 4'hd, 4'h4, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h5, 4'h0, 4'hf, 4'h4, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'h1, 4'hd, 4'hd, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'hc, 4'h0, 4'hd };
assign dw_0[660] = dw_0_660[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_661 = { 4'hf, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'hd, 4'h4, 4'h4, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'h7, 4'h1, 4'h0, 4'hc, 4'h5, 4'h0, 4'h4, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h4, 4'h3, 4'h3, 4'h4, 4'h0, 4'h5, 4'h1, 4'hc, 4'h0, 4'h3, 4'h0, 4'h1, 4'hd, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'hc, 4'h1, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1 };
assign dw_0[661] = dw_0_661[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_662 = { 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'hd, 4'h4, 4'h4, 4'h4, 4'h3, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'hd, 4'h3, 4'h3, 4'h4, 4'h5, 4'hf, 4'h3, 4'h4, 4'h0, 4'h4, 4'h1, 4'hf, 4'h4, 4'h3, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1 };
assign dw_0[662] = dw_0_662[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_663 = { 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'h4, 4'h7, 4'h3, 4'hc, 4'hd, 4'h1, 4'hd, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'h1, 4'h4, 4'hc, 4'h7, 4'h0, 4'h4, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'hd, 4'h3, 4'h3, 4'h0, 4'h7, 4'h3, 4'h3, 4'h4, 4'h0, 4'h5, 4'h1, 4'hf, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'h3, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1 };
assign dw_0[663] = dw_0_663[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_664 = { 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'hd, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h7, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h7, 4'h0, 4'h1, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0, 4'h5, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'hd, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h3, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'hd };
assign dw_0[664] = dw_0_664[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_665 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h7, 4'h3, 4'hc, 4'hd, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h7, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h7, 4'h3, 4'hc, 4'h3, 4'h3, 4'h4, 4'h4, 4'hf, 4'h7, 4'h0, 4'h0, 4'h5, 4'h1, 4'hf, 4'h4, 4'h0, 4'h1, 4'h4, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'hf, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1 };
assign dw_0[665] = dw_0_665[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_666 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h4, 4'hd, 4'h4, 4'h0, 4'h7, 4'h3, 4'hc, 4'hd, 4'h0, 4'hd, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h7, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'h3, 4'h3, 4'hd, 4'h3, 4'h3, 4'h4, 4'h5, 4'h3, 4'h4, 4'h4, 4'h0, 4'h5, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'hd, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd };
assign dw_0[666] = dw_0_666[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_667 = { 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'hf, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'h1, 4'hd, 4'h0, 4'h1, 4'h1, 4'h7, 4'h0, 4'h7, 4'hc, 4'h4, 4'h0, 4'h5, 4'h5, 4'h7, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h5, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[667] = dw_0_667[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_668 = { 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'hf, 4'h3, 4'h7, 4'h3, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'hc, 4'h4, 4'hc, 4'h1, 4'h7, 4'h0, 4'h3, 4'hd, 4'h4, 4'h0, 4'h5, 4'h1, 4'h4, 4'hc, 4'hc, 4'h3, 4'h1, 4'hf, 4'h4, 4'h3, 4'hf, 4'h4, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h1, 4'hc, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[668] = dw_0_668[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_669 = { 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hd, 4'h3, 4'h4, 4'h3, 4'h3, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'h1, 4'h4, 4'hd, 4'h5, 4'h7, 4'h0, 4'h3, 4'hc, 4'h4, 4'h0, 4'h4, 4'h1, 4'h4, 4'h1, 4'hd, 4'h3, 4'h1, 4'hc, 4'h5, 4'h0, 4'h0, 4'hc, 4'h4, 4'h5, 4'h0, 4'h7, 4'h0, 4'h0, 4'hc, 4'h1, 4'hd, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h1, 4'hc, 4'hd, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[669] = dw_0_669[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_670 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'hd, 4'h4, 4'h4, 4'h3, 4'h4, 4'hc, 4'h1, 4'h1, 4'hd, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h4, 4'hc, 4'hf, 4'hc, 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'hd, 4'h3, 4'h1, 4'hc, 4'h1, 4'h7, 4'h3, 4'hc, 4'h4, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'hf, 4'h1, 4'hd, 4'h1, 4'h0, 4'h4, 4'h0, 4'h4, 4'h7, 4'h1, 4'hd, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3 };
assign dw_0[670] = dw_0_670[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_671 = { 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'hd, 4'h4, 4'h0, 4'hf, 4'h3, 4'hc, 4'hd, 4'hc, 4'hd, 4'h1, 4'h1, 4'hd, 4'h1, 4'hc, 4'h1, 4'h4, 4'h0, 4'hf, 4'h3, 4'h7, 4'h0, 4'h4, 4'hd, 4'h4, 4'h0, 4'hc, 4'h3, 4'h1, 4'h0, 4'h5, 4'h7, 4'h0, 4'hc, 4'h4, 4'h1, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h1, 4'h3, 4'h1, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf };
assign dw_0[671] = dw_0_671[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_672 = { 4'h1, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h7, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h5, 4'hd, 4'h1, 4'hf, 4'h5, 4'h7, 4'h3, 4'h0, 4'h4, 4'h3, 4'hc, 4'h0, 4'h7, 4'h0, 4'hf, 4'h4, 4'hd, 4'h1, 4'h4, 4'hc, 4'h0, 4'h1, 4'h3, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'h5, 4'h1, 4'hc, 4'hf };
assign dw_0[672] = dw_0_672[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_673 = { 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h7, 4'h0, 4'h4, 4'h1, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h4, 4'h5, 4'hd, 4'h3, 4'hf, 4'h1, 4'h3, 4'h3, 4'h3, 4'h0, 4'hf, 4'hc, 4'h3, 4'h7, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc };
assign dw_0[673] = dw_0_673[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_674 = { 4'hd, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h3, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'h5, 4'h4, 4'h5, 4'hd, 4'h0, 4'hf, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc };
assign dw_0[674] = dw_0_674[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_675 = { 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h1, 4'h4, 4'h5, 4'hd, 4'h0, 4'h3, 4'h5, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc };
assign dw_0[675] = dw_0_675[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_676 = { 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'h1, 4'hd, 4'h3, 4'h0, 4'h5, 4'h0, 4'h5, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h4, 4'h5, 4'hc, 4'h0, 4'hf, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h4, 4'h3, 4'h0, 4'h3, 4'h1, 4'h1, 4'h3, 4'h5, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'hc, 4'hc };
assign dw_0[676] = dw_0_676[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_677 = { 4'h1, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h7, 4'h4, 4'h4, 4'h5, 4'hd, 4'h0, 4'hf, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc };
assign dw_0[677] = dw_0_677[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_678 = { 4'h1, 4'h7, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h4, 4'h0, 4'h5, 4'h0, 4'h5, 4'h3, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'h7, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hd, 4'h4, 4'h0, 4'h4, 4'h5, 4'hd, 4'h0, 4'hf, 4'h5, 4'h7, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'hd, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'hc };
assign dw_0[678] = dw_0_678[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_679 = { 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'hd, 4'h3, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hd, 4'h3, 4'h0, 4'h4, 4'h5, 4'hd, 4'h3, 4'hc, 4'h1, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h1, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc };
assign dw_0[679] = dw_0_679[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_680 = { 4'h1, 4'h7, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'h7, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h7, 4'h5, 4'h0, 4'h5, 4'hd, 4'h3, 4'hf, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h7, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h3, 4'hc, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[680] = dw_0_680[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_681 = { 4'h1, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'hc, 4'h1, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h7, 4'h5, 4'h4, 4'h5, 4'hd, 4'h3, 4'h3, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h7, 4'h0, 4'hf, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc };
assign dw_0[681] = dw_0_681[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_682 = { 4'h1, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'h5, 4'h0, 4'h3, 4'h1, 4'hc, 4'h0, 4'h0, 4'hf, 4'h1, 4'h1, 4'hc, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h5, 4'h4, 4'h5, 4'hd, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc };
assign dw_0[682] = dw_0_682[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_683 = { 4'h1, 4'h7, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h5, 4'h1, 4'h4, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'hc, 4'h3, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'hc };
assign dw_0[683] = dw_0_683[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_684 = { 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'hd, 4'hd, 4'h7, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h4, 4'hd, 4'h0, 4'hf, 4'h1, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h7, 4'h0, 4'h3, 4'h1, 4'h1, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc };
assign dw_0[684] = dw_0_684[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_685 = { 4'h1, 4'h7, 4'h4, 4'h3, 4'h0, 4'h1, 4'h1, 4'h7, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h4, 4'h4, 4'hd, 4'h3, 4'h3, 4'h1, 4'h3, 4'h3, 4'h3, 4'h0, 4'h7, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'hc, 4'h1, 4'h0, 4'h5, 4'hf, 4'h0, 4'h3, 4'hf, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc };
assign dw_0[685] = dw_0_685[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_686 = { 4'h1, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'hd, 4'h0, 4'hf, 4'h1, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'h3, 4'h4, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc };
assign dw_0[686] = dw_0_686[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_687 = { 4'h1, 4'h7, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h5, 4'hd, 4'h4, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h7, 4'h4, 4'h4, 4'h4, 4'hc, 4'h0, 4'hf, 4'h5, 4'h3, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'h0, 4'hf, 4'h0, 4'h1, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'hc };
assign dw_0[687] = dw_0_687[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_688 = { 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h7, 4'h5, 4'hf, 4'h1, 4'hf, 4'h7, 4'hf, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h4, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hd, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h3, 4'h7, 4'h1, 4'h7, 4'h5, 4'h0, 4'h1, 4'h4, 4'h3, 4'h1, 4'h0, 4'h1, 4'h7, 4'h7, 4'h1, 4'hf, 4'hf, 4'h0, 4'h1, 4'hf, 4'h0, 4'hf, 4'hf, 4'h1, 4'h0, 4'h0, 4'h7, 4'h0, 4'h1 };
assign dw_0[688] = dw_0_688[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_689 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h3, 4'hc, 4'h3, 4'h7, 4'hf, 4'h0, 4'h1, 4'h0, 4'h4, 4'hf, 4'h0, 4'hc, 4'h3, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'h7, 4'h3, 4'h3, 4'h3, 4'h5, 4'h0, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h3, 4'h1, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'hf, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h5 };
assign dw_0[689] = dw_0_689[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_690 = { 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h3, 4'h4, 4'hf, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h5, 4'h0, 4'h0, 4'h3, 4'h7, 4'h3, 4'hc, 4'h0, 4'h4, 4'hc, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'hf, 4'hf, 4'h0, 4'h1, 4'hc, 4'hc, 4'hf, 4'hf, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0 };
assign dw_0[690] = dw_0_690[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_691 = { 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h3, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h1, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h1, 4'hc, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h3, 4'h1, 4'hf, 4'hf, 4'h0, 4'h1, 4'hc, 4'hc, 4'hc, 4'hc, 4'hc, 4'h0, 4'h1, 4'h3, 4'h0, 4'h4 };
assign dw_0[691] = dw_0_691[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_692 = { 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'hf, 4'h3, 4'hf, 4'h0, 4'h1, 4'hd, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h3, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h0, 4'h7, 4'h0, 4'hf, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h7, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'hc, 4'h7 };
assign dw_0[692] = dw_0_692[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_693 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'h1, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h4, 4'hf, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'hd, 4'h4, 4'h3, 4'hd, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h1, 4'h0, 4'h1, 4'h3, 4'hc, 4'h4 };
assign dw_0[693] = dw_0_693[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_694 = { 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'h4, 4'hc, 4'h3, 4'h4, 4'h0, 4'h4, 4'hd, 4'h0, 4'h1, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h5, 4'hc, 4'hd, 4'h0, 4'hd, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h7, 4'h0, 4'h1, 4'hf, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3 };
assign dw_0[694] = dw_0_694[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_695 = { 4'h4, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'h1, 4'h0, 4'h5, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h3, 4'h5, 4'h0, 4'hf, 4'h7, 4'h5, 4'h0, 4'hd, 4'h0, 4'h1, 4'h4, 4'h1, 4'h5, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0 };
assign dw_0[695] = dw_0_695[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_696 = { 4'h7, 4'h7, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'h3, 4'hf, 4'hf, 4'hc, 4'h1, 4'hc, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h5, 4'h4, 4'h1, 4'h0, 4'h7, 4'h1, 4'h3, 4'h0, 4'h4, 4'h1, 4'h1, 4'h4, 4'hd, 4'h7, 4'h0, 4'hd, 4'h0, 4'hd, 4'h4, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h1, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3 };
assign dw_0[696] = dw_0_696[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_697 = { 4'h7, 4'h7, 4'hc, 4'h1, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'h1, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h4, 4'h7, 4'h4, 4'hc, 4'h1, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'h1, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h1, 4'h7, 4'h0, 4'hd, 4'h0, 4'hd, 4'h7, 4'h7, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3 };
assign dw_0[697] = dw_0_697[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_698 = { 4'h0, 4'h7, 4'h0, 4'h1, 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'h1, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'hf, 4'h1, 4'hc, 4'h4, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd, 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'hc, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h3, 4'h1, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0 };
assign dw_0[698] = dw_0_698[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_699 = { 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h7, 4'h4, 4'h3, 4'h1, 4'hf, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'h4, 4'h1, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h7, 4'h3, 4'h1, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0 };
assign dw_0[699] = dw_0_699[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_700 = { 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h5, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h7, 4'h4, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'hd, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0 };
assign dw_0[700] = dw_0_700[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_701 = { 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h7, 4'h4, 4'hf, 4'h0, 4'hf, 4'h0, 4'hf, 4'hc, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h7, 4'h4, 4'h3, 4'h3, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0 };
assign dw_0[701] = dw_0_701[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_702 = { 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h3, 4'h4, 4'hc, 4'h0, 4'hf, 4'h7, 4'hf, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h7, 4'h4, 4'h3, 4'hc, 4'h3, 4'h5, 4'h3, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h7, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'h1, 4'hf, 4'hc, 4'hf, 4'hf, 4'hd, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0 };
assign dw_0[702] = dw_0_702[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_703 = { 4'h3, 4'h3, 4'h4, 4'h1, 4'h0, 4'hf, 4'h4, 4'hf, 4'h5, 4'hf, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'h1, 4'hf, 4'h1, 4'h4, 4'h4, 4'hf, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'hd, 4'hc, 4'h1, 4'h3, 4'hc, 4'h4, 4'h3, 4'h7, 4'h7, 4'h0, 4'h7, 4'h5, 4'h0, 4'h1, 4'h5, 4'h3, 4'h0, 4'h1, 4'hc, 4'h4, 4'h7, 4'hc, 4'hf, 4'hf, 4'h0, 4'h1, 4'hf, 4'h0, 4'hc, 4'hf, 4'hd, 4'h0, 4'h4, 4'h7, 4'h0, 4'h1 };
assign dw_0[703] = dw_0_703[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_704 = { 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h1, 4'h4, 4'h5, 4'hc, 4'hc, 4'h4, 4'h3, 4'hc, 4'h7, 4'h5, 4'hd, 4'h3, 4'h3, 4'h0, 4'hf, 4'h4, 4'hc, 4'hf, 4'h0, 4'h5, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'hf, 4'h1, 4'h1, 4'hc, 4'h7, 4'hd, 4'h0, 4'hd, 4'hc, 4'h7, 4'h0, 4'h3, 4'hc, 4'h4, 4'hc, 4'h0, 4'h5, 4'h3, 4'h0, 4'hc, 4'hd, 4'h4, 4'h0, 4'h3, 4'hc, 4'h5, 4'h5, 4'h3, 4'h1, 4'h0, 4'h3, 4'hc, 4'h4, 4'h5 };
assign dw_0[704] = dw_0_704[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_705 = { 4'hd, 4'h5, 4'h4, 4'h1, 4'h0, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h7, 4'h1, 4'h5, 4'h1, 4'h1, 4'h1, 4'h0, 4'h4, 4'hc, 4'hc, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'hf, 4'h5, 4'h5, 4'h3, 4'h3, 4'h5, 4'h0, 4'hd, 4'h0, 4'h7, 4'h4, 4'h3, 4'hc, 4'h0, 4'hd, 4'h0, 4'h1, 4'hf, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h4, 4'h5 };
assign dw_0[705] = dw_0_705[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_706 = { 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h1, 4'h5, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'hc, 4'hc, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h1, 4'hf, 4'h5, 4'h5, 4'h7, 4'h3, 4'h5, 4'h0, 4'h1, 4'h4, 4'h3, 4'h0, 4'hf, 4'hc, 4'h1, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h4, 4'h4 };
assign dw_0[706] = dw_0_706[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_707 = { 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc, 4'h7, 4'h1, 4'h5, 4'h1, 4'h0, 4'h1, 4'h3, 4'h5, 4'hc, 4'hc, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h7, 4'h5, 4'hf, 4'h4, 4'h4, 4'hc, 4'h3, 4'h5, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hf, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4 };
assign dw_0[707] = dw_0_707[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_708 = { 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h1, 4'hc, 4'h4, 4'h4, 4'h7, 4'hc, 4'h0, 4'hc, 4'h7, 4'h1, 4'h5, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'hd, 4'hc, 4'h4, 4'h0, 4'h4, 4'h1, 4'hf, 4'h5, 4'h5, 4'h7, 4'h0, 4'h5, 4'h0, 4'h1, 4'h4, 4'hf, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h7, 4'h0, 4'h3, 4'h4, 4'h4, 4'h5, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h4, 4'h7 };
assign dw_0[708] = dw_0_708[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_709 = { 4'hc, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h3, 4'hd, 4'hc, 4'hc, 4'h4, 4'hd, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hd, 4'h1, 4'h4, 4'h0, 4'h4, 4'h1, 4'hf, 4'h5, 4'h5, 4'h0, 4'h1, 4'h5, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'h1, 4'hd, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'hd, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h0, 4'hd, 4'h0, 4'hf, 4'hf, 4'h4, 4'h4 };
assign dw_0[709] = dw_0_709[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_710 = { 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h5, 4'h3, 4'h3, 4'hd, 4'hc, 4'hc, 4'h4, 4'hd, 4'h5, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h3, 4'h4, 4'h5, 4'h0, 4'h1, 4'h5, 4'h3, 4'h1, 4'h1, 4'h3, 4'h0, 4'hf, 4'hf, 4'h1, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'h5, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'hf, 4'h3, 4'h4, 4'h7 };
assign dw_0[710] = dw_0_710[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_711 = { 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'h5, 4'h0, 4'h3, 4'hc, 4'hc, 4'hc, 4'h7, 4'h1, 4'h1, 4'h4, 4'h0, 4'h5, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'hd, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'hf, 4'h5, 4'h5, 4'h7, 4'h1, 4'h1, 4'h0, 4'h1, 4'h1, 4'hf, 4'h4, 4'hf, 4'hf, 4'h5, 4'hd, 4'h0, 4'hc, 4'h3, 4'h3, 4'h7, 4'h0, 4'h4, 4'h0, 4'h3, 4'h5, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h4, 4'h7 };
assign dw_0[711] = dw_0_711[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_712 = { 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'hf, 4'hc, 4'h3, 4'hc, 4'h4, 4'hd, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'hc, 4'h0, 4'hd, 4'h1, 4'h4, 4'h0, 4'h3, 4'h5, 4'hf, 4'h5, 4'h0, 4'h7, 4'h1, 4'h5, 4'h3, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h1, 4'hd, 4'h0, 4'h5, 4'hc, 4'h0, 4'h3, 4'hc, 4'h4, 4'h0, 4'h3, 4'h5, 4'h0, 4'h5, 4'hd, 4'hd, 4'h0, 4'hc, 4'h0, 4'h4, 4'h7 };
assign dw_0[712] = dw_0_712[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_713 = { 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h7, 4'hd, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'hc, 4'h4, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'hf, 4'h5, 4'h4, 4'h4, 4'h1, 4'h1, 4'h0, 4'h1, 4'h3, 4'h3, 4'h4, 4'hf, 4'h3, 4'h5, 4'h3, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h7, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4 };
assign dw_0[713] = dw_0_713[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_714 = { 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h5, 4'h0, 4'h0, 4'hd, 4'h1, 4'hd, 4'h7, 4'hd, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hd, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'hf, 4'h5, 4'h4, 4'h3, 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'hf, 4'h4, 4'hf, 4'hf, 4'h5, 4'h0, 4'h0, 4'hd, 4'h3, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'h4, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7 };
assign dw_0[714] = dw_0_714[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_715 = { 4'hc, 4'h5, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'h3, 4'h0, 4'h7, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hd, 4'h1, 4'h4, 4'h0, 4'h4, 4'h4, 4'hf, 4'h5, 4'h5, 4'h3, 4'h0, 4'h4, 4'h3, 4'hd, 4'h3, 4'h3, 4'h0, 4'hf, 4'hc, 4'h5, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h7, 4'h5, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4 };
assign dw_0[715] = dw_0_715[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_716 = { 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hc, 4'hc, 4'hc, 4'h1, 4'h0, 4'h4, 4'h4, 4'h4, 4'h4, 4'hf, 4'h5, 4'h5, 4'h3, 4'h0, 4'h5, 4'h3, 4'hd, 4'h0, 4'h3, 4'h4, 4'hf, 4'hc, 4'h1, 4'hc, 4'h0, 4'hd, 4'hc, 4'h0, 4'h3, 4'h1, 4'h7, 4'h0, 4'h3, 4'h5, 4'h4, 4'h5, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4 };
assign dw_0[716] = dw_0_716[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_717 = { 4'hc, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'hd, 4'hc, 4'h0, 4'h0, 4'hc, 4'h7, 4'h4, 4'h5, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'hc, 4'hc, 4'hc, 4'h1, 4'h1, 4'h4, 4'h0, 4'h5, 4'h1, 4'hf, 4'h0, 4'h5, 4'h3, 4'h3, 4'h5, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'h5, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h4, 4'h4 };
assign dw_0[717] = dw_0_717[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_718 = { 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h5, 4'h5, 4'h1, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h1, 4'h4, 4'hc, 4'h4, 4'h4, 4'hf, 4'h5, 4'h5, 4'h3, 4'hf, 4'h5, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'hf, 4'hd, 4'h1, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5 };
assign dw_0[718] = dw_0_718[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_719 = { 4'hc, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'hc, 4'hf, 4'h4, 4'hc, 4'hc, 4'h4, 4'h1, 4'h5, 4'h3, 4'h3, 4'h0, 4'h3, 4'h5, 4'hc, 4'hc, 4'h0, 4'h5, 4'h1, 4'h5, 4'h0, 4'h4, 4'h4, 4'hf, 4'h5, 4'h5, 4'h3, 4'h3, 4'h1, 4'h3, 4'hd, 4'hd, 4'h7, 4'h0, 4'h3, 4'h1, 4'h1, 4'hc, 4'h0, 4'h1, 4'hf, 4'h3, 4'h0, 4'hd, 4'h7, 4'h0, 4'hf, 4'h1, 4'h4, 4'h5, 4'h3, 4'h1, 4'h0, 4'h0, 4'hf, 4'h4, 4'h5 };
assign dw_0[719] = dw_0_719[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_720 = { 4'h1, 4'h0, 4'h4, 4'h3, 4'h0, 4'hf, 4'hd, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h1, 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h4, 4'h4, 4'h7, 4'h4, 4'h1, 4'hd, 4'h1, 4'hc, 4'h5, 4'h3, 4'h5, 4'h0, 4'h4, 4'h4, 4'h0, 4'h7, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h7, 4'h7, 4'h1, 4'h0, 4'h4, 4'h5, 4'h3, 4'h1, 4'hc, 4'h4, 4'h0, 4'h1, 4'h3, 4'h0, 4'hd };
assign dw_0[720] = dw_0_720[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_721 = { 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'hd, 4'h0, 4'hc, 4'h1, 4'hf, 4'h0, 4'h0, 4'hc, 4'h1, 4'h1, 4'h1, 4'h0, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h4, 4'h1, 4'h3, 4'h1, 4'h1, 4'hc, 4'h1, 4'hd, 4'h5, 4'h3, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h7, 4'h0, 4'h7, 4'h3, 4'hd, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'h5, 4'h7, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd };
assign dw_0[721] = dw_0_721[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_722 = { 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h7, 4'h1, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h4, 4'h1, 4'h7, 4'h1, 4'h1, 4'hc, 4'h1, 4'h0, 4'h1, 4'h3, 4'h5, 4'h0, 4'h0, 4'h1, 4'hc, 4'h7, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h7, 4'h1, 4'h0, 4'h3, 4'h4, 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc };
assign dw_0[722] = dw_0_722[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_723 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hd, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h5, 4'h1, 4'h1, 4'h1, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h7, 4'h1, 4'h0, 4'h3, 4'h5, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd };
assign dw_0[723] = dw_0_723[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_724 = { 4'hc, 4'h1, 4'h4, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'h3, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'h7, 4'h1, 4'h1, 4'hc, 4'h0, 4'hc, 4'h5, 4'h3, 4'h4, 4'h3, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h7, 4'h1, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'hd };
assign dw_0[724] = dw_0_724[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_725 = { 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'hd, 4'hc, 4'h1, 4'h1, 4'h4, 4'h0, 4'hc, 4'hf, 4'h0, 4'h5, 4'h1, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'hc, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'h5, 4'h4, 4'h7, 4'h1, 4'h1, 4'h1, 4'h3, 4'hc, 4'h1, 4'h3, 4'h5, 4'h5, 4'h0, 4'h5, 4'h0, 4'h7, 4'hc, 4'h3, 4'h3, 4'hc, 4'h1, 4'h0, 4'h7, 4'h1, 4'h0, 4'h3, 4'h5, 4'h3, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd };
assign dw_0[725] = dw_0_725[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_726 = { 4'hc, 4'h1, 4'h4, 4'h3, 4'h0, 4'h3, 4'hc, 4'h1, 4'hc, 4'h4, 4'h4, 4'h0, 4'hc, 4'hc, 4'h1, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hd, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h7, 4'h5, 4'h5, 4'h1, 4'h3, 4'hc, 4'h5, 4'h3, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h5, 4'h7, 4'h4, 4'h0, 4'h3, 4'h1, 4'h3, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd };
assign dw_0[726] = dw_0_726[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_727 = { 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'hc, 4'hf, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'hc, 4'h3, 4'h3, 4'h4, 4'h0, 4'h4, 4'hc, 4'h3, 4'h1, 4'h5, 4'h0, 4'h3, 4'hc, 4'h5, 4'h3, 4'h4, 4'h4, 4'hc, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h1, 4'hf, 4'h1, 4'h0, 4'h0, 4'hc, 4'hc, 4'hd };
assign dw_0[727] = dw_0_727[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_728 = { 4'h0, 4'hd, 4'h4, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h1, 4'h5, 4'h1, 4'h1, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h4, 4'h0, 4'h5, 4'h4, 4'h4, 4'h1, 4'h5, 4'h1, 4'h3, 4'h0, 4'h1, 4'h3, 4'h5, 4'h5, 4'h0, 4'h4, 4'h1, 4'h4, 4'h3, 4'h0, 4'hf, 4'hc, 4'hd, 4'h0, 4'h7, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1, 4'hf, 4'h1, 4'h0, 4'h0, 4'hc, 4'hc, 4'hd };
assign dw_0[728] = dw_0_728[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_729 = { 4'h3, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h5, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'h7, 4'h3, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h1, 4'h0, 4'hc, 4'h4, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'hd };
assign dw_0[729] = dw_0_729[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_730 = { 4'h0, 4'h1, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'hf, 4'h1, 4'h5, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h7, 4'h3, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'h7, 4'h5, 4'h0, 4'h0, 4'h1, 4'hf, 4'hd, 4'hc, 4'h1, 4'h0, 4'h4, 4'hc, 4'h0, 4'hd };
assign dw_0[730] = dw_0_730[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_731 = { 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'hf, 4'h0, 4'h4, 4'h1, 4'h0, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h7, 4'h3, 4'h4, 4'h0, 4'h4, 4'h0, 4'h7, 4'h1, 4'h5, 4'h1, 4'h3, 4'hc, 4'h4, 4'h3, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h4, 4'h7, 4'h5, 4'h0, 4'h3, 4'h0, 4'hf, 4'h1, 4'hc, 4'h1, 4'h0, 4'h1, 4'hc, 4'h0, 4'hd };
assign dw_0[731] = dw_0_731[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_732 = { 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h5, 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h3, 4'h4, 4'h0, 4'h5, 4'h0, 4'h3, 4'h1, 4'h5, 4'h1, 4'h0, 4'h1, 4'h4, 4'h3, 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4, 4'hc, 4'hd, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hd };
assign dw_0[732] = dw_0_732[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_733 = { 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'hc, 4'h1, 4'h4, 4'h1, 4'h0, 4'h7, 4'h3, 4'hd, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h5, 4'h1, 4'h3, 4'h1, 4'h1, 4'h1, 4'h1, 4'hc, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h3, 4'h3, 4'hc, 4'hd, 4'h4, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hd };
assign dw_0[733] = dw_0_733[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_734 = { 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'hd, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h1, 4'hf, 4'h1, 4'h3, 4'h1, 4'hc, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h7, 4'h5, 4'h0, 4'h0, 4'h5, 4'h3, 4'hd, 4'h1, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc };
assign dw_0[734] = dw_0_734[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_735 = { 4'h0, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'hd, 4'hc, 4'h4, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h1, 4'h1, 4'h0, 4'hc, 4'h3, 4'h1, 4'h0, 4'hc, 4'h4, 4'h3, 4'h3, 4'h4, 4'h0, 4'h5, 4'h1, 4'h3, 4'h1, 4'h5, 4'hc, 4'h1, 4'hf, 4'h4, 4'h7, 4'h5, 4'hd, 4'hc, 4'h0, 4'h1, 4'h7, 4'h3, 4'h3, 4'h4, 4'h0, 4'h1, 4'h5, 4'h7, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'hd, 4'hd, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc };
assign dw_0[735] = dw_0_735[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_736 = { 4'hc, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h7, 4'h3, 4'h1, 4'h0, 4'hf, 4'hc, 4'h0, 4'h1, 4'h0, 4'h4, 4'h7, 4'h3, 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'hd, 4'hf, 4'hc, 4'hc, 4'h0, 4'hc, 4'hf, 4'h3, 4'hc, 4'hd, 4'h3, 4'hd, 4'hc, 4'h0, 4'hf, 4'h3, 4'h5, 4'h0, 4'h3, 4'hc, 4'hc, 4'h4, 4'h0, 4'h7, 4'h0, 4'hf, 4'hf, 4'h4, 4'h0 };
assign dw_0[736] = dw_0_736[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_737 = { 4'hc, 4'h5, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h5, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h7, 4'h7, 4'h0, 4'h4, 4'h5, 4'h4, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h3, 4'hd, 4'h3, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4 };
assign dw_0[737] = dw_0_737[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_738 = { 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h1, 4'h1, 4'h4, 4'h0, 4'h7, 4'h3, 4'h1, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'h5, 4'h4, 4'h0, 4'h1, 4'hf, 4'hc, 4'hc, 4'h1, 4'h0, 4'hc, 4'h3, 4'hc, 4'h1, 4'h3, 4'hd, 4'hc, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3 };
assign dw_0[738] = dw_0_738[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_739 = { 4'hc, 4'h4, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h1, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h3, 4'h1, 4'h0, 4'hd, 4'hf, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4 };
assign dw_0[739] = dw_0_739[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_740 = { 4'hf, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h1, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h3, 4'h1, 4'h0, 4'h1, 4'hc, 4'h0, 4'h3, 4'hc, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0 };
assign dw_0[740] = dw_0_740[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_741 = { 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h1, 4'hc, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'hd, 4'h5, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h1, 4'h0, 4'hd, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'hc, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0 };
assign dw_0[741] = dw_0_741[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_742 = { 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h3, 4'h1, 4'h4, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hd, 4'h4, 4'h5, 4'h4, 4'h0, 4'h3, 4'hc, 4'hc, 4'hc, 4'h1, 4'hc, 4'hc, 4'h0, 4'h3, 4'h1, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4 };
assign dw_0[742] = dw_0_742[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_743 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h7, 4'h3, 4'h1, 4'h4, 4'hf, 4'hc, 4'hc, 4'hd, 4'h0, 4'h0, 4'hf, 4'h4, 4'h3, 4'h4, 4'h5, 4'h5, 4'h0, 4'h1, 4'hf, 4'hc, 4'h1, 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'h5, 4'h0, 4'h0, 4'hd, 4'hf, 4'h1, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4 };
assign dw_0[743] = dw_0_743[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_744 = { 4'h1, 4'h4, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h1, 4'h4, 4'hf, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'h7, 4'h4, 4'h3, 4'h1, 4'h5, 4'hc, 4'h1, 4'hc, 4'hc, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h3, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0 };
assign dw_0[744] = dw_0_744[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_745 = { 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h7, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h4, 4'h0, 4'h5, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h1, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0 };
assign dw_0[745] = dw_0_745[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_746 = { 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h4, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h4, 4'h5, 4'h5, 4'h0, 4'h1, 4'hc, 4'hc, 4'h1, 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'h3, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h4 };
assign dw_0[746] = dw_0_746[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_747 = { 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'hd, 4'h0, 4'hd, 4'hc, 4'h0, 4'hc, 4'hc, 4'h1, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0 };
assign dw_0[747] = dw_0_747[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_748 = { 4'h0, 4'h5, 4'hc, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h1, 4'h4, 4'h1, 4'h0, 4'h7, 4'h3, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h7, 4'h1, 4'h4, 4'h1, 4'h4, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'hc, 4'h5, 4'h0, 4'h3, 4'hd, 4'hf, 4'h5, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4 };
assign dw_0[748] = dw_0_748[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_749 = { 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'h1, 4'hd, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h7, 4'h3, 4'h0, 4'h4, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h1, 4'hc, 4'hc, 4'hd, 4'hc, 4'hc, 4'hc, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'h3, 4'hc, 4'h3, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0 };
assign dw_0[749] = dw_0_749[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_750 = { 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'h3, 4'h1, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hd, 4'hc, 4'hf, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'hd, 4'h4, 4'h4 };
assign dw_0[750] = dw_0_750[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_751 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h1, 4'h4, 4'hf, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h4, 4'h4, 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'hd, 4'h4, 4'h3, 4'h1, 4'h0, 4'hd, 4'hc, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd, 4'h0, 4'h1, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h4 };
assign dw_0[751] = dw_0_751[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_752 = { 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'hf, 4'h5, 4'hc, 4'h4, 4'hc, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'hf, 4'h1, 4'h0, 4'h4, 4'h0, 4'h4, 4'h4, 4'h7, 4'h0, 4'h3, 4'hd, 4'h4, 4'hc, 4'h3, 4'h5, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'hc, 4'hf, 4'h3, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hd, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h1, 4'hf, 4'h0, 4'h1 };
assign dw_0[752] = dw_0_752[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_753 = { 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h1, 4'h0, 4'hc, 4'h3, 4'h4, 4'h0, 4'h4, 4'h1, 4'h7, 4'h4, 4'h5, 4'h5, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'hf, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'hd, 4'h3, 4'h0, 4'h0, 4'h1, 4'hf, 4'hc, 4'h1 };
assign dw_0[753] = dw_0_753[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_754 = { 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h4, 4'hd, 4'hc, 4'h3, 4'h0, 4'h5, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h7, 4'h0, 4'h0, 4'h5, 4'h4, 4'hc, 4'h3, 4'h0, 4'h1, 4'h4, 4'h1, 4'h7, 4'h0, 4'h4, 4'h5, 4'hd, 4'hf, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h1 };
assign dw_0[754] = dw_0_754[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_755 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hd, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h1, 4'h0, 4'hc, 4'h1, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'hc, 4'hf, 4'h5, 4'h4, 4'hc, 4'h0, 4'h3, 4'h1, 4'h4, 4'h1, 4'h3, 4'h0, 4'h5, 4'h1, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'hf, 4'h1, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[755] = dw_0_755[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_756 = { 4'h3, 4'hc, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hd, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h1, 4'hc, 4'h0, 4'hf, 4'hc, 4'h5, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h7, 4'h0, 4'hf, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h4, 4'h4, 4'h1, 4'hc, 4'h0, 4'h4, 4'hf, 4'hf, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0 };
assign dw_0[756] = dw_0_756[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_757 = { 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hd, 4'hc, 4'h1, 4'h0, 4'h5, 4'h0, 4'h1, 4'h1, 4'h0, 4'hf, 4'hc, 4'h5, 4'h4, 4'hf, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h4, 4'hc, 4'h1, 4'h1, 4'h1, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h7, 4'hf, 4'h3, 4'h1, 4'h4, 4'h5, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0 };
assign dw_0[757] = dw_0_757[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_758 = { 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hd, 4'hc, 4'h0, 4'hc, 4'h5, 4'h0, 4'h1, 4'hc, 4'h0, 4'hf, 4'h0, 4'h5, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'hd, 4'hc, 4'h0, 4'h1, 4'h7, 4'h1, 4'hd, 4'h3, 4'h5, 4'hc, 4'hc, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'h1, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0 };
assign dw_0[758] = dw_0_758[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_759 = { 4'h3, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'hf, 4'hd, 4'hc, 4'hc, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'hc, 4'h4, 4'h4, 4'hf, 4'h3, 4'h0, 4'h0, 4'h7, 4'h3, 4'hc, 4'h1, 4'h4, 4'hd, 4'h1, 4'h0, 4'h0, 4'h7, 4'h1, 4'hf, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h5, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0 };
assign dw_0[759] = dw_0_759[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_760 = { 4'h0, 4'hd, 4'hc, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'hc, 4'hd, 4'h0, 4'h5, 4'h1, 4'h1, 4'hc, 4'h1, 4'hf, 4'hc, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'h5, 4'h0, 4'h1, 4'h4, 4'hc, 4'h1, 4'h0, 4'hd, 4'h4, 4'h1, 4'hf, 4'h4, 4'h0, 4'h3, 4'hd, 4'h3, 4'h0, 4'h7, 4'hc, 4'hc, 4'h5, 4'h7, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3 };
assign dw_0[760] = dw_0_760[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_761 = { 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'hc, 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'h5, 4'hd, 4'h1, 4'hc, 4'h1, 4'h4, 4'h1, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3 };
assign dw_0[761] = dw_0_761[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_762 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'hc, 4'h3, 4'h3, 4'h0, 4'hc, 4'hd, 4'hc, 4'h1, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'hc, 4'h1, 4'h5, 4'hc, 4'h1, 4'h3, 4'h1, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0 };
assign dw_0[762] = dw_0_762[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_763 = { 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'hf, 4'hd, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'hc, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'hc, 4'h1, 4'h4, 4'hc, 4'h1, 4'h0, 4'h1, 4'h4, 4'h1, 4'h3, 4'h4, 4'h4, 4'h0, 4'h1, 4'hf, 4'h3, 4'h0, 4'hc, 4'hf, 4'h5, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0 };
assign dw_0[763] = dw_0_763[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_764 = { 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hd, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h4, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'hc, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0 };
assign dw_0[764] = dw_0_764[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_765 = { 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'hc, 4'hf, 4'hc, 4'h3, 4'hd, 4'hc, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h1, 4'h4, 4'h3, 4'h3, 4'h4, 4'h0, 4'h5, 4'hc, 4'hc, 4'h1, 4'h5, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'hc, 4'h0, 4'h3, 4'h4, 4'hc, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1 };
assign dw_0[765] = dw_0_765[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_766 = { 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hd, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'hd, 4'h1, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h4, 4'hc, 4'hc, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h1, 4'h7, 4'h4, 4'h4, 4'h1, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1 };
assign dw_0[766] = dw_0_766[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_767 = { 4'h0, 4'hc, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h1, 4'hc, 4'h5, 4'h0, 4'h1, 4'hd, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'h5, 4'h5, 4'hd, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h1, 4'hf, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hd, 4'h3, 4'hc, 4'h3, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1 };
assign dw_0[767] = dw_0_767[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_768 = { 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'h7, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h7, 4'h7, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0 };
assign dw_0[768] = dw_0_768[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_769 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h1, 4'hc, 4'h0, 4'hc, 4'h1, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf };
assign dw_0[769] = dw_0_769[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_770 = { 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h4, 4'h0, 4'h5, 4'h0, 4'h3, 4'h7, 4'hd, 4'h1, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc, 4'h3 };
assign dw_0[770] = dw_0_770[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_771 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h1, 4'h7, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h5, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h1, 4'hc, 4'hf, 4'hd, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0 };
assign dw_0[771] = dw_0_771[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_772 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h1, 4'hc, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'hf };
assign dw_0[772] = dw_0_772[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_773 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'h4, 4'hc, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0 };
assign dw_0[773] = dw_0_773[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_774 = { 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'hf, 4'h1, 4'hc, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h5, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0 };
assign dw_0[774] = dw_0_774[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_775 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h5, 4'h0, 4'h3, 4'hd, 4'h0, 4'hf, 4'h0, 4'hc, 4'hf, 4'h1, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0 };
assign dw_0[775] = dw_0_775[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_776 = { 4'hc, 4'hc, 4'h4, 4'h3, 4'h0, 4'h1, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'hc, 4'hf, 4'h1, 4'hc, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h0 };
assign dw_0[776] = dw_0_776[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_777 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'hc, 4'h3, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0 };
assign dw_0[777] = dw_0_777[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_778 = { 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[778] = dw_0_778[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_779 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'hd, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0 };
assign dw_0[779] = dw_0_779[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_780 = { 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h7, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'h1, 4'h1, 4'h0, 4'h0, 4'h7, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'hf, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'h7, 4'hc, 4'hc, 4'h1, 4'h1, 4'h1, 4'h0, 4'h3, 4'h3, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[780] = dw_0_780[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_781 = { 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd, 4'hc, 4'h4, 4'hf, 4'h4, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'hd, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'hc, 4'h1, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3 };
assign dw_0[781] = dw_0_781[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_782 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h5, 4'hc, 4'h3, 4'hd, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h1, 4'hc, 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'h7, 4'hc, 4'hc, 4'h5, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h3, 4'h7, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'hc, 4'h3 };
assign dw_0[782] = dw_0_782[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_783 = { 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'hf, 4'h7, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h3, 4'hc, 4'h3, 4'hc, 4'h1, 4'hf, 4'hf, 4'hd, 4'hc, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h7, 4'h4, 4'h1, 4'h0, 4'h1, 4'hc, 4'hc, 4'hc };
assign dw_0[783] = dw_0_783[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_784 = { 4'h0, 4'h7, 4'h4, 4'h3, 4'h0, 4'h7, 4'hd, 4'h3, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'hd, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'hd, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'h3, 4'h7, 4'h4, 4'h0, 4'h0, 4'h5, 4'h3, 4'hf, 4'h4, 4'h3, 4'h3, 4'h1, 4'h4, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h7, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'hf };
assign dw_0[784] = dw_0_784[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_785 = { 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'hf, 4'h7, 4'h4, 4'hc, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h1, 4'h4, 4'h3, 4'h7, 4'h3, 4'h1, 4'h0, 4'hc, 4'hd, 4'hd, 4'h7, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc };
assign dw_0[785] = dw_0_785[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_786 = { 4'h3, 4'h7, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h1, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h1, 4'h4, 4'h5, 4'h7, 4'h7, 4'h1, 4'h0, 4'hf, 4'hd, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h3, 4'h3, 4'h3, 4'h0, 4'hd, 4'h1, 4'hc, 4'hc };
assign dw_0[786] = dw_0_786[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_787 = { 4'h0, 4'h7, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'hc, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'hd, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'h1, 4'h4, 4'h4, 4'h7, 4'h3, 4'h1, 4'h0, 4'hc, 4'hd, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'h1, 4'hc, 4'hc };
assign dw_0[787] = dw_0_787[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_788 = { 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h4, 4'hc, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h7, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'hf, 4'h0, 4'h3, 4'hf, 4'h1, 4'h4, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'hd, 4'hd, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hf, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc };
assign dw_0[788] = dw_0_788[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_789 = { 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h7, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'hf, 4'h1, 4'h3, 4'hf, 4'h1, 4'h4, 4'h7, 4'h7, 4'h3, 4'h0, 4'h0, 4'hd, 4'hd, 4'hd, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'hc, 4'hc };
assign dw_0[789] = dw_0_789[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_790 = { 4'h1, 4'h7, 4'h4, 4'h3, 4'h0, 4'h4, 4'h1, 4'h3, 4'h0, 4'h4, 4'hf, 4'h5, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h4, 4'hc, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h7, 4'h7, 4'h3, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'hf, 4'hf, 4'h1, 4'h4, 4'h5, 4'h4, 4'h3, 4'h5, 4'h0, 4'hd, 4'hc, 4'h0, 4'h3, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0 };
assign dw_0[790] = dw_0_790[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_791 = { 4'h3, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h7, 4'h0, 4'hc, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h5, 4'h4, 4'h3, 4'h1, 4'h0, 4'h1, 4'hd, 4'h0, 4'h3, 4'h7, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'hc, 4'hc };
assign dw_0[791] = dw_0_791[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_792 = { 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'hf, 4'h4, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hd, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h7, 4'h0, 4'h3, 4'h4, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'h0, 4'h4, 4'h5, 4'h4, 4'h3, 4'h5, 4'h0, 4'hc, 4'hd, 4'h1, 4'h0, 4'h7, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'hf };
assign dw_0[792] = dw_0_792[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_793 = { 4'h0, 4'h7, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h5, 4'h4, 4'h1, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'h4, 4'hc, 4'hc, 4'h7, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'h4, 4'h4, 4'h7, 4'h3, 4'h4, 4'h0, 4'hd, 4'hd, 4'hc, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'hd, 4'h0, 4'hc };
assign dw_0[793] = dw_0_793[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_794 = { 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h5, 4'h4, 4'h1, 4'h0, 4'hf, 4'h0, 4'h3, 4'hf, 4'h3, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'h7, 4'h0, 4'hf, 4'hd, 4'h3, 4'hf, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h5, 4'h0, 4'hd, 4'hd, 4'h0, 4'h7, 4'h4, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[794] = dw_0_794[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_795 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'hd, 4'h3, 4'hf, 4'h4, 4'h4, 4'h4, 4'h0, 4'h7, 4'h0, 4'h0, 4'hc, 4'hd, 4'h1, 4'h4, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'hd, 4'h0, 4'h0 };
assign dw_0[795] = dw_0_795[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_796 = { 4'h0, 4'h7, 4'h4, 4'h3, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc, 4'h5, 4'h4, 4'hd, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h7, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'h1, 4'h4, 4'h4, 4'h3, 4'h3, 4'h1, 4'h0, 4'hd, 4'hd, 4'hd, 4'h3, 4'h4, 4'h5, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc };
assign dw_0[796] = dw_0_796[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_797 = { 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h7, 4'h3, 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'h1, 4'h4, 4'h4, 4'h7, 4'h7, 4'h1, 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[797] = dw_0_797[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_798 = { 4'h1, 4'h7, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h1, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'hd, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h3, 4'hf, 4'h1, 4'h4, 4'h4, 4'h4, 4'h3, 4'h1, 4'h0, 4'hd, 4'hd, 4'h0, 4'h3, 4'h7, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0 };
assign dw_0[798] = dw_0_798[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_799 = { 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h1, 4'h0, 4'hd, 4'h0, 4'hc, 4'h3, 4'h3, 4'h3, 4'h3, 4'h5, 4'h0, 4'h1, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h7, 4'h7, 4'h0, 4'hc, 4'h7, 4'h3, 4'hc, 4'h4, 4'h3, 4'h3, 4'h4, 4'h4, 4'h4, 4'h0, 4'h3, 4'h5, 4'h1, 4'hd, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'hd, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc };
assign dw_0[799] = dw_0_799[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_800 = { 4'hd, 4'hd, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'hf, 4'h0, 4'h4, 4'hf, 4'h0, 4'h1, 4'h0, 4'h4, 4'h3, 4'h3, 4'h4, 4'h3, 4'h1, 4'h1, 4'h7, 4'h4, 4'h4, 4'h1, 4'hc, 4'hc, 4'h5, 4'h7, 4'h5, 4'hd, 4'hc, 4'h1, 4'h7, 4'hc, 4'hf, 4'h4, 4'hf, 4'h4, 4'h0, 4'h5, 4'h7, 4'hd, 4'hc, 4'h3, 4'h5, 4'hf, 4'h0, 4'h5, 4'hc, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h3, 4'h5, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0 };
assign dw_0[800] = dw_0_800[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_801 = { 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'h4, 4'hf, 4'h0, 4'h4, 4'h4, 4'h4, 4'hd, 4'h1, 4'hc, 4'h3, 4'h5, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'hc, 4'h4, 4'h0, 4'h5, 4'h4, 4'hc, 4'h0, 4'h5, 4'h3, 4'h7, 4'h3, 4'h1, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'hd, 4'hc, 4'h0, 4'h1, 4'hf, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h7, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h3, 4'hc, 4'h3 };
assign dw_0[801] = dw_0_801[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_802 = { 4'h1, 4'hd, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'hf, 4'h3, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'hd, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'hc, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'h1, 4'h3, 4'h1, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'h5, 4'hd, 4'hd, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3 };
assign dw_0[802] = dw_0_802[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_803 = { 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h5, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'h4, 4'h1, 4'h0, 4'h5, 4'h0, 4'h3, 4'h3, 4'h0, 4'h7, 4'hd, 4'hc, 4'h5, 4'h4, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h3, 4'h7, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'hc, 4'h3 };
assign dw_0[803] = dw_0_803[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_804 = { 4'hc, 4'h1, 4'hc, 4'h1, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'hf, 4'h0, 4'h5, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'hc, 4'h0, 4'h5, 4'h0, 4'h4, 4'hd, 4'hc, 4'h5, 4'h0, 4'h3, 4'hc, 4'hd, 4'h3, 4'h1, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'h4, 4'hf, 4'h0, 4'h1, 4'hd, 4'hd, 4'h0, 4'h3, 4'h3, 4'h4, 4'h7, 4'h0, 4'h1, 4'h0, 4'hf, 4'h3, 4'h0, 4'h3 };
assign dw_0[804] = dw_0_804[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_805 = { 4'h0, 4'h7, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'h5, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'hd, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'h1, 4'h4, 4'h3, 4'hc, 4'h0, 4'h3, 4'h1, 4'hc, 4'h1, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'h3, 4'h3, 4'h5, 4'h4, 4'hc, 4'h1, 4'h0, 4'hf, 4'h3, 4'h0, 4'h3 };
assign dw_0[805] = dw_0_805[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_806 = { 4'h1, 4'h0, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h0, 4'h4, 4'h3, 4'hd, 4'h0, 4'h0, 4'h4, 4'h5, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h4, 4'h3, 4'hc, 4'h0, 4'h7, 4'hd, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h7, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf };
assign dw_0[806] = dw_0_806[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_807 = { 4'hd, 4'h4, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'hc, 4'hf, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h1, 4'h0, 4'h4, 4'h4, 4'h1, 4'h1, 4'hc, 4'h0, 4'h1, 4'h1, 4'h4, 4'hf, 4'hd, 4'h1, 4'h4, 4'hf, 4'h0, 4'hd, 4'h3, 4'hd, 4'hc, 4'h1, 4'h0, 4'hd, 4'hc, 4'h0, 4'h1, 4'hf, 4'h0, 4'hc, 4'hc, 4'hd, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3 };
assign dw_0[807] = dw_0_807[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_808 = { 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'h5, 4'h3, 4'h1, 4'h5, 4'hc, 4'hf, 4'hf, 4'h0, 4'h4, 4'h7, 4'h4, 4'hd, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'h1, 4'h4, 4'h4, 4'hc, 4'hf, 4'h5, 4'h0, 4'h3, 4'hc, 4'hd, 4'h7, 4'h1, 4'hc, 4'h5, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'hd, 4'hc, 4'hd, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3 };
assign dw_0[808] = dw_0_808[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_809 = { 4'hc, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h3, 4'h1, 4'h5, 4'hc, 4'h3, 4'hf, 4'h0, 4'h5, 4'h4, 4'h4, 4'hd, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'h4, 4'h5, 4'h1, 4'hc, 4'h0, 4'h1, 4'h4, 4'h4, 4'hc, 4'hf, 4'h5, 4'h0, 4'h3, 4'hc, 4'h1, 4'h7, 4'h1, 4'hc, 4'h5, 4'h0, 4'h1, 4'hc, 4'h3, 4'hc, 4'hf, 4'h0, 4'h1, 4'h1, 4'hd, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3 };
assign dw_0[809] = dw_0_809[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_810 = { 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'h7, 4'h0, 4'h1, 4'h5, 4'h0, 4'hc, 4'hf, 4'h0, 4'h4, 4'h0, 4'h4, 4'hc, 4'h1, 4'h7, 4'h0, 4'h1, 4'h4, 4'h3, 4'h0, 4'h5, 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'h4, 4'hc, 4'h3, 4'h5, 4'h1, 4'h3, 4'h0, 4'h0, 4'h7, 4'h1, 4'hc, 4'h1, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hd, 4'hd, 4'h0, 4'h3, 4'h3, 4'h1, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7 };
assign dw_0[810] = dw_0_810[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_811 = { 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'h1, 4'h4, 4'hc, 4'hc, 4'hf, 4'h4, 4'h4, 4'h0, 4'h4, 4'hc, 4'h1, 4'h1, 4'h3, 4'hd, 4'h4, 4'h7, 4'h0, 4'h5, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h0, 4'h7, 4'h0, 4'hc, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3 };
assign dw_0[811] = dw_0_811[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_812 = { 4'hd, 4'hc, 4'hc, 4'h1, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h5, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'hf, 4'h1, 4'h4, 4'h4, 4'h0, 4'h5, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'hd, 4'h3, 4'h5, 4'h0, 4'hf, 4'h0, 4'hd, 4'h7, 4'h5, 4'hc, 4'h1, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'hd, 4'hd, 4'hc, 4'h0, 4'h3, 4'h4, 4'h4, 4'h3, 4'h0, 4'hd, 4'h0, 4'hf, 4'hf, 4'h0, 4'h3 };
assign dw_0[812] = dw_0_812[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_813 = { 4'hc, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'hf, 4'h4, 4'h5, 4'h1, 4'hc, 4'h0, 4'h0, 4'h5, 4'hc, 4'hc, 4'h3, 4'h5, 4'h0, 4'hf, 4'h3, 4'hd, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'hd, 4'hd, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h4, 4'h3 };
assign dw_0[813] = dw_0_813[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_814 = { 4'h1, 4'h1, 4'hc, 4'h1, 4'h0, 4'h7, 4'h3, 4'h1, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'hc, 4'h3, 4'hd, 4'h3, 4'h1, 4'h4, 4'h7, 4'h4, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'hf, 4'h5, 4'h3, 4'hf, 4'hc, 4'h1, 4'h3, 4'h5, 4'hc, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'hf, 4'h0, 4'hc, 4'h1, 4'hd, 4'h0, 4'h3, 4'hf, 4'h5, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0 };
assign dw_0[814] = dw_0_814[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_815 = { 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'h4, 4'h1, 4'h1, 4'hf, 4'hd, 4'h7, 4'hf, 4'h1, 4'h4, 4'h4, 4'h5, 4'hf, 4'h3, 4'h7, 4'h3, 4'h1, 4'h0, 4'h4, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'h5, 4'h4, 4'hf, 4'hf, 4'h4, 4'hc, 4'h4, 4'hc, 4'h5, 4'h7, 4'h1, 4'hc, 4'h3, 4'h1, 4'hf, 4'hc, 4'h1, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'h4, 4'h7, 4'h5, 4'h0, 4'h3, 4'hf, 4'h0, 4'h1 };
assign dw_0[815] = dw_0_815[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_816 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd, 4'h0, 4'hf, 4'h1, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h1, 4'h0, 4'h5, 4'h4, 4'h5, 4'hd, 4'h4, 4'hc, 4'h3, 4'h4, 4'h4, 4'h0, 4'hc, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'hf, 4'hc, 4'h1, 4'h3, 4'h0, 4'h1, 4'h5, 4'h0, 4'h3 };
assign dw_0[816] = dw_0_816[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_817 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'h1, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h3, 4'hd, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7 };
assign dw_0[817] = dw_0_817[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_818 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hc, 4'h7, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h4, 4'h1, 4'h4, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h7, 4'h4, 4'h0, 4'hc, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h3, 4'hf, 4'hc, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3 };
assign dw_0[818] = dw_0_818[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_819 = { 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'h5, 4'h0, 4'hf, 4'h4, 4'h4, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0 };
assign dw_0[819] = dw_0_819[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_820 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h1, 4'h1, 4'h0, 4'h5, 4'h4, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4 };
assign dw_0[820] = dw_0_820[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_821 = { 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h4, 4'h4, 4'h4, 4'h1, 4'h5, 4'h5, 4'h0, 4'hc, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4 };
assign dw_0[821] = dw_0_821[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_822 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h1, 4'h1, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h3, 4'h4, 4'h4, 4'h1, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0 };
assign dw_0[822] = dw_0_822[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_823 = { 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'hd, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h5, 4'h0, 4'h3, 4'h4, 4'h4, 4'h5, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h3, 4'h0, 4'h1, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h5 };
assign dw_0[823] = dw_0_823[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_824 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h4, 4'h4, 4'h5, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'hf, 4'h3, 4'h0, 4'h4, 4'h0, 4'h7, 4'h4, 4'h0, 4'h5, 4'h1, 4'h4, 4'h4, 4'h0, 4'hc, 4'h4, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'hf, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5 };
assign dw_0[824] = dw_0_824[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_825 = { 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'h1, 4'hd, 4'h0, 4'h1, 4'h5, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'h7, 4'h5, 4'h0, 4'h1, 4'h1, 4'h7, 4'h4, 4'h0, 4'hd, 4'h7, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1 };
assign dw_0[825] = dw_0_825[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_826 = { 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h3, 4'h3, 4'h5, 4'h0, 4'h3, 4'h4, 4'h4, 4'h5, 4'h1, 4'h7, 4'h4, 4'h0, 4'hc, 4'h7, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[826] = dw_0_826[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_827 = { 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'hc, 4'h7, 4'h0, 4'h0, 4'h4, 4'h1, 4'h3, 4'h4, 4'h4, 4'h1, 4'h1, 4'h4, 4'h4, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h1, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4 };
assign dw_0[827] = dw_0_827[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_828 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h1, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h1, 4'hc, 4'h5, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'hc, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1 };
assign dw_0[828] = dw_0_828[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_829 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'hc, 4'h1, 4'hf, 4'h0, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'h5, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0 };
assign dw_0[829] = dw_0_829[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_830 = { 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h3, 4'h1, 4'h4, 4'h3, 4'h1, 4'h0, 4'h5, 4'h4, 4'h4, 4'hc, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'hc, 4'h1, 4'h3, 4'h0, 4'h5, 4'h1, 4'h0, 4'h4 };
assign dw_0[830] = dw_0_830[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_831 = { 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'hc, 4'h4, 4'hc, 4'h0, 4'h0, 4'hd, 4'h1, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h1, 4'h0, 4'h3, 4'h1, 4'h0, 4'h5, 4'h4, 4'h4, 4'hc, 4'h4, 4'hf, 4'h3, 4'h7, 4'h4, 4'h0, 4'hc, 4'h7, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'hc, 4'hd, 4'hd, 4'h3, 4'h0, 4'h5, 4'h5, 4'h0, 4'h3 };
assign dw_0[831] = dw_0_831[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_832 = { 4'h1, 4'h3, 4'hc, 4'h1, 4'h0, 4'h3, 4'h3, 4'h5, 4'hc, 4'h4, 4'h0, 4'h7, 4'hc, 4'hf, 4'h0, 4'hd, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'hf, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h1, 4'hf, 4'h1, 4'hf, 4'h3, 4'h7, 4'h1, 4'h1, 4'hc, 4'h3, 4'h0, 4'h7, 4'h0, 4'hf, 4'hc, 4'h3, 4'h4, 4'h1, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'h5, 4'h7, 4'h1, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc };
assign dw_0[832] = dw_0_832[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_833 = { 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h7, 4'h3, 4'h0, 4'hc, 4'h4, 4'h1, 4'h7, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h4, 4'h0, 4'hc, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'h7, 4'hc, 4'hf, 4'hf, 4'hf, 4'h7, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h7, 4'h0, 4'h4, 4'h0, 4'h7, 4'h4, 4'h0, 4'hc };
assign dw_0[833] = dw_0_833[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_834 = { 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h4, 4'hf, 4'h3, 4'h4, 4'h4, 4'hd, 4'h3, 4'h1, 4'hf, 4'hc, 4'hc, 4'h4, 4'h0, 4'hc, 4'h5, 4'h1, 4'hc, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'h1, 4'hc, 4'h3, 4'h3, 4'hf, 4'hc, 4'hf, 4'hc, 4'hf, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'hc, 4'h5, 4'h7, 4'hc, 4'h5, 4'h0, 4'h7, 4'h0, 4'hc, 4'hf };
assign dw_0[834] = dw_0_834[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_835 = { 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h7, 4'h0, 4'h4, 4'hd, 4'h3, 4'hd, 4'hf, 4'hd, 4'hc, 4'h4, 4'h3, 4'hf, 4'h5, 4'h5, 4'hd, 4'hf, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'hf, 4'h3, 4'h0, 4'h1, 4'hc, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'hd, 4'h3, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'hc, 4'h5, 4'h4, 4'h0, 4'h5, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0 };
assign dw_0[835] = dw_0_835[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_836 = { 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h7, 4'h1, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h4, 4'h3, 4'h3, 4'h5, 4'h1, 4'hd, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h1, 4'hc, 4'h3, 4'hc, 4'h7, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0, 4'h7, 4'hc, 4'h5, 4'h7, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'hc, 4'hf };
assign dw_0[836] = dw_0_836[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_837 = { 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'hf, 4'h4, 4'h3, 4'h4, 4'h1, 4'h3, 4'h0, 4'hf, 4'hd, 4'hd, 4'h4, 4'h3, 4'h3, 4'h4, 4'h1, 4'hc, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h1, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'h7, 4'hc, 4'hf, 4'hc, 4'h3, 4'h4, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h7, 4'h1, 4'hc, 4'hc };
assign dw_0[837] = dw_0_837[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_838 = { 4'h4, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h4, 4'h1, 4'h3, 4'h0, 4'hf, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'hf, 4'h4, 4'hf, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h4, 4'hc, 4'h3, 4'hc, 4'h3, 4'hc, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'hc, 4'h5, 4'h0, 4'h0, 4'hc, 4'h1, 4'h7, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc };
assign dw_0[838] = dw_0_838[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_839 = { 4'h5, 4'h4, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'h3, 4'h1, 4'hf, 4'h0, 4'hd, 4'h7, 4'h3, 4'h0, 4'h0, 4'h5, 4'hc, 4'hf, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h5, 4'hf, 4'h0, 4'h4, 4'h0, 4'h1, 4'hc, 4'hf, 4'hc, 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'h3, 4'h1, 4'hd, 4'hf, 4'h0, 4'h5, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'h7, 4'hc, 4'h5, 4'h0, 4'h7, 4'h0, 4'h0, 4'hf };
assign dw_0[839] = dw_0_839[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_840 = { 4'h4, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'hd, 4'h3, 4'h1, 4'h3, 4'hd, 4'h1, 4'h3, 4'h3, 4'h0, 4'h1, 4'h5, 4'hd, 4'h3, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'hc, 4'h3, 4'h1, 4'h3, 4'h4, 4'hf, 4'h0, 4'h5, 4'hc, 4'hf, 4'hc, 4'h3, 4'hc, 4'hf, 4'hc, 4'hf, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h7, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'hc, 4'hf };
assign dw_0[840] = dw_0_840[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_841 = { 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h3, 4'h1, 4'h4, 4'h7, 4'h1, 4'h3, 4'h0, 4'hf, 4'hc, 4'hd, 4'h3, 4'h0, 4'hf, 4'h5, 4'h0, 4'hd, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'hf, 4'h5, 4'hf, 4'h3, 4'h7, 4'h0, 4'h1, 4'hc, 4'h3, 4'h3, 4'h7, 4'h0, 4'hf, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hf, 4'h1, 4'h0, 4'h0, 4'hf, 4'h1, 4'h7, 4'h1, 4'h0, 4'h0, 4'h7, 4'h3, 4'h0, 4'hf };
assign dw_0[841] = dw_0_841[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_842 = { 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h1, 4'h3, 4'h4, 4'hd, 4'h4, 4'h1, 4'hf, 4'hc, 4'hd, 4'h7, 4'h0, 4'hf, 4'h5, 4'h0, 4'hd, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h5, 4'hf, 4'h7, 4'h4, 4'h0, 4'h1, 4'hd, 4'hf, 4'hc, 4'h7, 4'h0, 4'hf, 4'hc, 4'hf, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h5, 4'h7, 4'hc, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'hf };
assign dw_0[842] = dw_0_842[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_843 = { 4'h5, 4'h1, 4'h0, 4'h1, 4'h0, 4'h7, 4'h3, 4'h1, 4'h0, 4'h4, 4'h1, 4'h7, 4'h1, 4'hf, 4'hc, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'hf, 4'h0, 4'hf, 4'h3, 4'h7, 4'h4, 4'hd, 4'h3, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc, 4'hf, 4'hc, 4'h7, 4'hc, 4'hf, 4'hc, 4'h3, 4'h4, 4'h0, 4'h4, 4'hd, 4'h0, 4'hc, 4'hf, 4'h4, 4'h0, 4'hf, 4'h1, 4'h5, 4'h4, 4'hf, 4'h1, 4'h0, 4'h7, 4'hc, 4'h0, 4'hc };
assign dw_0[843] = dw_0_843[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_844 = { 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc, 4'h7, 4'h3, 4'h4, 4'h1, 4'h4, 4'h4, 4'h3, 4'hd, 4'hd, 4'h4, 4'h3, 4'hf, 4'h4, 4'h0, 4'hc, 4'hf, 4'h4, 4'hf, 4'h3, 4'h3, 4'h4, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3, 4'h5, 4'hc, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hc, 4'hf, 4'h4, 4'h0, 4'h4, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h4, 4'hf, 4'h5, 4'h7, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3 };
assign dw_0[844] = dw_0_844[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_845 = { 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'hd, 4'h7, 4'hc, 4'hf, 4'hd, 4'hc, 4'h0, 4'h0, 4'hc, 4'h5, 4'h1, 4'hc, 4'hf, 4'h0, 4'hf, 4'hf, 4'h3, 4'h4, 4'hd, 4'h3, 4'hd, 4'h3, 4'h0, 4'h7, 4'h3, 4'h4, 4'hc, 4'hf, 4'hf, 4'h0, 4'hc, 4'hf, 4'hd, 4'h3, 4'h1, 4'h1, 4'h0, 4'hc, 4'h0, 4'h1, 4'hf, 4'h5, 4'h0, 4'h4, 4'hd, 4'h5, 4'h4, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'hc, 4'hf };
assign dw_0[845] = dw_0_845[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_846 = { 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'hc, 4'hf, 4'h3, 4'h5, 4'h7, 4'h1, 4'h3, 4'h0, 4'hf, 4'h0, 4'hc, 4'h5, 4'h1, 4'hc, 4'h5, 4'h1, 4'hc, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h4, 4'h7, 4'h0, 4'h4, 4'hd, 4'hf, 4'h7, 4'h3, 4'hc, 4'hf, 4'hc, 4'hf, 4'h4, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'hc, 4'h5, 4'h7, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf };
assign dw_0[846] = dw_0_846[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_847 = { 4'h4, 4'h3, 4'hc, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'hd, 4'h4, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'hd, 4'h4, 4'h1, 4'hc, 4'h0, 4'h1, 4'hd, 4'hf, 4'h0, 4'hf, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h5, 4'hc, 4'h3, 4'h4, 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h7, 4'hd, 4'h1, 4'h0, 4'h3, 4'h4, 4'h0, 4'hf };
assign dw_0[847] = dw_0_847[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_848 = { 4'h4, 4'hd, 4'h4, 4'h3, 4'h0, 4'h3, 4'hf, 4'hc, 4'hd, 4'h7, 4'h3, 4'h5, 4'hd, 4'hd, 4'h0, 4'hd, 4'h3, 4'h3, 4'hd, 4'h0, 4'h4, 4'h5, 4'h4, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h1, 4'hc, 4'h4, 4'hf, 4'hd, 4'hd, 4'h7, 4'hf, 4'h4, 4'h7, 4'h7, 4'h3, 4'h4, 4'h1, 4'hd, 4'hf, 4'h7, 4'h1, 4'h7, 4'h5, 4'h5, 4'h1, 4'h3, 4'h5, 4'h0, 4'h1, 4'h4, 4'h4, 4'hc, 4'h0, 4'h3, 4'h0, 4'h5, 4'h5, 4'hc, 4'hc };
assign dw_0[848] = dw_0_848[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_849 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h1, 4'h0, 4'hc, 4'h4, 4'hc, 4'h1, 4'h0, 4'hd, 4'hc, 4'hc, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'hc, 4'h7, 4'hc, 4'h3, 4'h4, 4'h4, 4'hf, 4'h3, 4'h7, 4'h0, 4'h7, 4'h1, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc };
assign dw_0[849] = dw_0_849[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_850 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h1, 4'h1, 4'hd, 4'h5, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc, 4'h0, 4'hd, 4'h4, 4'hf, 4'h0, 4'h7, 4'hf, 4'h7, 4'h4, 4'h4, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h7, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc, 4'hc };
assign dw_0[850] = dw_0_850[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_851 = { 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h1, 4'h1, 4'hd, 4'h0, 4'hc, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'hf, 4'h4, 4'h3, 4'h0, 4'hd, 4'h0, 4'hf, 4'h0, 4'h7, 4'hf, 4'h7, 4'h0, 4'h4, 4'h3, 4'hf, 4'h3, 4'h0, 4'h7, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc };
assign dw_0[851] = dw_0_851[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_852 = { 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h1, 4'h4, 4'h3, 4'h1, 4'h0, 4'hd, 4'h0, 4'hc, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'hf, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hd, 4'hc, 4'h0, 4'h7, 4'hd, 4'h7, 4'h0, 4'h3, 4'h4, 4'h5, 4'h3, 4'h0, 4'h7, 4'h0, 4'h4, 4'h1, 4'hc, 4'h3, 4'h7, 4'hc, 4'h4, 4'h0, 4'h3, 4'h1, 4'h1, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc };
assign dw_0[852] = dw_0_852[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_853 = { 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h7, 4'h5, 4'h3, 4'hc, 4'hd, 4'h0, 4'hd, 4'hc, 4'hc, 4'h1, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hd, 4'h3, 4'h7, 4'h4, 4'h5, 4'hc, 4'h3, 4'h5, 4'h0, 4'h7, 4'h0, 4'hf, 4'h4, 4'h5, 4'h0, 4'hc, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'hd, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc };
assign dw_0[853] = dw_0_853[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_854 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h5, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hc, 4'h7, 4'hf, 4'h3, 4'h4, 4'h5, 4'h0, 4'hf, 4'h3, 4'h0, 4'h7, 4'h0, 4'h1, 4'h1, 4'h7, 4'h1, 4'h0, 4'h0, 4'h7, 4'h5, 4'hc, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'hc, 4'hc };
assign dw_0[854] = dw_0_854[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_855 = { 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hd, 4'h4, 4'h0, 4'h3, 4'h1, 4'h4, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'h0, 4'hc, 4'hd, 4'h3, 4'h3, 4'hc, 4'h4, 4'h3, 4'h7, 4'h4, 4'h5, 4'h0, 4'hc, 4'hf, 4'h0, 4'hc, 4'hd, 4'hc, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc };
assign dw_0[855] = dw_0_855[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_856 = { 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'hf, 4'hc, 4'hd, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'hd, 4'hc, 4'hc, 4'h0, 4'h3, 4'hd, 4'h5, 4'h0, 4'hc, 4'h5, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h7, 4'h3, 4'h0, 4'hd, 4'h0, 4'hf, 4'hc, 4'h4, 4'hf, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0 };
assign dw_0[856] = dw_0_856[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_857 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h5, 4'h0, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'h1, 4'h1, 4'hd, 4'h1, 4'h0, 4'h0, 4'h5, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'hd, 4'h0, 4'h7, 4'hc, 4'h4, 4'h3, 4'h3, 4'h4, 4'h4, 4'h0, 4'hf, 4'h7, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc };
assign dw_0[857] = dw_0_857[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_858 = { 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'hf, 4'hd, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'hd, 4'h0, 4'hc, 4'h1, 4'h0, 4'hc, 4'h1, 4'h1, 4'h1, 4'h1, 4'hc, 4'h3, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h7, 4'h4, 4'h7, 4'h4, 4'h4, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'hc };
assign dw_0[858] = dw_0_858[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_859 = { 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'hd, 4'h0, 4'hc, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'hc, 4'hd, 4'h0, 4'h3, 4'h0, 4'h7, 4'h3, 4'h7, 4'h4, 4'h4, 4'hc, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc };
assign dw_0[859] = dw_0_859[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_860 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hd, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h4, 4'h0, 4'hc, 4'hd, 4'h0, 4'hf, 4'hc, 4'h7, 4'hf, 4'h7, 4'h4, 4'h4, 4'hf, 4'h3, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc };
assign dw_0[860] = dw_0_860[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_861 = { 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h3, 4'hd, 4'h1, 4'h0, 4'hc, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hd, 4'h4, 4'h0, 4'h0, 4'hd, 4'h4, 4'hc, 4'h1, 4'h7, 4'hc, 4'h7, 4'h4, 4'h4, 4'hc, 4'h3, 4'h3, 4'h0, 4'h7, 4'h1, 4'h1, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h3, 4'h0, 4'hc };
assign dw_0[861] = dw_0_861[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_862 = { 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0, 4'h3, 4'hd, 4'h1, 4'h5, 4'h0, 4'h5, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h4, 4'h0, 4'h7, 4'hd, 4'h3, 4'hf, 4'hc, 4'h4, 4'hc, 4'h7, 4'h4, 4'h5, 4'hc, 4'hc, 4'h3, 4'h0, 4'h7, 4'h1, 4'h0, 4'hd, 4'h3, 4'h1, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc };
assign dw_0[862] = dw_0_862[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_863 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'hd, 4'hd, 4'hf, 4'h3, 4'h3, 4'hc, 4'h3, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h3, 4'h5, 4'h3, 4'h4, 4'hd, 4'h7, 4'hc, 4'h0, 4'h7, 4'hf, 4'h7, 4'h4, 4'h4, 4'hc, 4'hf, 4'h3, 4'h1, 4'h0, 4'h5, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0, 4'h1, 4'hc, 4'hd, 4'hd, 4'h4, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc };
assign dw_0[863] = dw_0_863[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_864 = { 4'h3, 4'h3, 4'hc, 4'h1, 4'h0, 4'h7, 4'h4, 4'hf, 4'h5, 4'hc, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h1, 4'h4, 4'h4, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h1, 4'h4, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0 };
assign dw_0[864] = dw_0_864[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_865 = { 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'h7, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h5, 4'h0, 4'h3, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h7, 4'h5, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h7, 4'h0, 4'h1 };
assign dw_0[865] = dw_0_865[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_866 = { 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hd, 4'hd, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h1, 4'hd, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1 };
assign dw_0[866] = dw_0_866[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_867 = { 4'h3, 4'h3, 4'hc, 4'h1, 4'h0, 4'h7, 4'h7, 4'hc, 4'hd, 4'h4, 4'h3, 4'h0, 4'hc, 4'h1, 4'h4, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'hd, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc };
assign dw_0[867] = dw_0_867[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_868 = { 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h7, 4'h0, 4'h7, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'h0, 4'h1, 4'h3, 4'h0, 4'hc };
assign dw_0[868] = dw_0_868[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_869 = { 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'h4, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h7, 4'hc, 4'h1, 4'h0, 4'h4, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0 };
assign dw_0[869] = dw_0_869[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_870 = { 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h4, 4'h3, 4'h0, 4'h1, 4'h1, 4'h4, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h7, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0 };
assign dw_0[870] = dw_0_870[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_871 = { 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0, 4'hc, 4'hd, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h7, 4'h0, 4'h4, 4'h4, 4'hc, 4'h4, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'h7, 4'h0, 4'h1, 4'h0, 4'h4, 4'hc };
assign dw_0[871] = dw_0_871[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_872 = { 4'h3, 4'h4, 4'hc, 4'h0, 4'h0, 4'h7, 4'h4, 4'hc, 4'hd, 4'h7, 4'hc, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3 };
assign dw_0[872] = dw_0_872[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_873 = { 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'hd, 4'h4, 4'h0, 4'h3, 4'hc, 4'hd, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h4, 4'h4, 4'h4, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'hd, 4'h0, 4'h3, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0 };
assign dw_0[873] = dw_0_873[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_874 = { 4'h7, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'h1, 4'h1, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h7, 4'hc, 4'h7, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3 };
assign dw_0[874] = dw_0_874[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_875 = { 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h7, 4'h0, 4'hd, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h4, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'hf, 4'hc, 4'h3, 4'hc, 4'h1, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3 };
assign dw_0[875] = dw_0_875[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_876 = { 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h5, 4'h0, 4'h4, 4'h0, 4'h4, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3 };
assign dw_0[876] = dw_0_876[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_877 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h7, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h5, 4'h5, 4'hf, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf };
assign dw_0[877] = dw_0_877[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_878 = { 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'hd, 4'hd, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h7, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3 };
assign dw_0[878] = dw_0_878[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_879 = { 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h7, 4'h4, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'hf, 4'hd, 4'h4, 4'hc, 4'h3, 4'h1, 4'hc, 4'h0, 4'h3, 4'h4, 4'hf, 4'hc, 4'h7, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'hf, 4'h5, 4'h4, 4'hf, 4'h4, 4'h3, 4'h4, 4'hc, 4'hd, 4'hf, 4'hc, 4'h0, 4'h1, 4'h4, 4'h7, 4'hf, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'h0, 4'hf, 4'hd, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3 };
assign dw_0[879] = dw_0_879[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_880 = { 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hd, 4'h3, 4'h4, 4'h5, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h7, 4'hf, 4'h0, 4'h4, 4'h3, 4'hc, 4'h1, 4'h5, 4'hc, 4'h0, 4'h3, 4'h7, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'hf, 4'hc, 4'hc, 4'hf, 4'h1, 4'hc, 4'hd, 4'h4, 4'h1, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h1, 4'h1, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h7, 4'h7, 4'h0, 4'hf, 4'h1, 4'h0, 4'h4 };
assign dw_0[880] = dw_0_880[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_881 = { 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'hd, 4'h1, 4'h7, 4'h0, 4'h0, 4'h3, 4'h7, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h5, 4'h4, 4'h3, 4'hc, 4'hd, 4'h1, 4'hc, 4'h0, 4'h3, 4'h4, 4'h5, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'hc, 4'hd, 4'hf, 4'h0, 4'hc, 4'hc, 4'h7, 4'h0, 4'h1, 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h1, 4'h3, 4'h4, 4'h3, 4'h0, 4'hf, 4'hd, 4'h0, 4'h4 };
assign dw_0[881] = dw_0_881[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_882 = { 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h3, 4'h1, 4'h4, 4'h3, 4'hc, 4'hd, 4'h4, 4'hc, 4'h0, 4'h3, 4'h4, 4'h5, 4'h3, 4'h0, 4'h4, 4'h0, 4'h3, 4'hf, 4'hd, 4'hf, 4'h1, 4'hc, 4'hd, 4'h3, 4'h1, 4'h1, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h3, 4'h4, 4'h3, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0 };
assign dw_0[882] = dw_0_882[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_883 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h1, 4'hc, 4'h0, 4'h3, 4'h7, 4'h3, 4'h1, 4'h4, 4'h3, 4'hc, 4'h1, 4'h5, 4'h0, 4'h0, 4'hf, 4'h4, 4'h5, 4'h7, 4'h0, 4'h5, 4'h0, 4'hc, 4'hc, 4'hd, 4'h3, 4'h1, 4'hc, 4'h1, 4'h4, 4'h0, 4'h5, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'h1, 4'h0, 4'h7 };
assign dw_0[883] = dw_0_883[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_884 = { 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h5, 4'h4, 4'h1, 4'h3, 4'h0, 4'h3, 4'h7, 4'h3, 4'h1, 4'h0, 4'h3, 4'hc, 4'h1, 4'h1, 4'h0, 4'h0, 4'hf, 4'h4, 4'h5, 4'h3, 4'hf, 4'h5, 4'h0, 4'h3, 4'h0, 4'hd, 4'hf, 4'h0, 4'hc, 4'hd, 4'h4, 4'h0, 4'h5, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'h1, 4'hc, 4'h3, 4'h4, 4'h3, 4'h0, 4'hf, 4'h1, 4'h4, 4'h0 };
assign dw_0[884] = dw_0_884[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_885 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h4, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'h3, 4'h7, 4'h3, 4'h0, 4'h4, 4'h7, 4'hc, 4'h1, 4'h5, 4'hc, 4'h0, 4'hf, 4'h4, 4'h5, 4'h3, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'hd, 4'hf, 4'h1, 4'hc, 4'hd, 4'h3, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'h4, 4'h3, 4'h0, 4'hf, 4'h1, 4'h4, 4'h0 };
assign dw_0[885] = dw_0_885[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_886 = { 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'hd, 4'hf, 4'h4, 4'h4, 4'h4, 4'hc, 4'hf, 4'h0, 4'h3, 4'h7, 4'h3, 4'h0, 4'h4, 4'h3, 4'hc, 4'h1, 4'h1, 4'h0, 4'h0, 4'hf, 4'h4, 4'h1, 4'h3, 4'hc, 4'h5, 4'h0, 4'h3, 4'h0, 4'hd, 4'h3, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'hd, 4'hf, 4'h1, 4'hf, 4'h1, 4'h1, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'hf, 4'h1, 4'h0, 4'h4 };
assign dw_0[886] = dw_0_886[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_887 = { 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'h4, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h7, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'h5, 4'h0, 4'h0, 4'hf, 4'h4, 4'h5, 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'hc, 4'hd, 4'h3, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0 };
assign dw_0[887] = dw_0_887[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_888 = { 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'hc, 4'h3, 4'h4, 4'h5, 4'h4, 4'h0, 4'hf, 4'h0, 4'h3, 4'h7, 4'h3, 4'h0, 4'h4, 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h4, 4'h5, 4'h3, 4'hf, 4'h5, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h4, 4'h5, 4'h0, 4'h1, 4'hc, 4'h0, 4'hc, 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h1, 4'h4, 4'h0 };
assign dw_0[888] = dw_0_888[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_889 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'hf, 4'h1, 4'h3, 4'h7, 4'h5, 4'h4, 4'h0, 4'hf, 4'h0, 4'h3, 4'h7, 4'h3, 4'h1, 4'h4, 4'h4, 4'hc, 4'h1, 4'h5, 4'h3, 4'h0, 4'hf, 4'h4, 4'h1, 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'hf, 4'h1, 4'h0, 4'h0, 4'h3, 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h1, 4'h1, 4'h0, 4'h3, 4'h1, 4'hc, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'h1, 4'h4, 4'h3 };
assign dw_0[889] = dw_0_889[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_890 = { 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h5, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h7, 4'h3, 4'h1, 4'h4, 4'h0, 4'hc, 4'h1, 4'h1, 4'h0, 4'h0, 4'hf, 4'h7, 4'h4, 4'h7, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'hd, 4'hf, 4'h1, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'hf, 4'h1, 4'h0, 4'h3 };
assign dw_0[890] = dw_0_890[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_891 = { 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h5, 4'hc, 4'h0, 4'h0, 4'h3, 4'h7, 4'h3, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h5, 4'h3, 4'hc, 4'h5, 4'h0, 4'h0, 4'hc, 4'hd, 4'hf, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'hf, 4'h0, 4'hc, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'h1, 4'h4, 4'h7 };
assign dw_0[891] = dw_0_891[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_892 = { 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'hc, 4'hf, 4'h7, 4'h5, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h7, 4'h3, 4'h1, 4'h4, 4'h3, 4'hc, 4'h1, 4'h1, 4'hc, 4'h0, 4'hf, 4'h4, 4'h5, 4'h3, 4'hc, 4'h4, 4'h0, 4'hc, 4'hc, 4'hd, 4'hf, 4'h5, 4'hc, 4'hd, 4'h4, 4'h0, 4'h1, 4'h0, 4'hd, 4'hc, 4'h0, 4'hf, 4'h1, 4'h1, 4'h0, 4'h3, 4'hd, 4'hc, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0 };
assign dw_0[892] = dw_0_892[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_893 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'h0, 4'h4, 4'h3, 4'hc, 4'h1, 4'h5, 4'hc, 4'h0, 4'hf, 4'h4, 4'h5, 4'h3, 4'hc, 4'h5, 4'h0, 4'h0, 4'hf, 4'hd, 4'hc, 4'h0, 4'hc, 4'hd, 4'h0, 4'h1, 4'h1, 4'h0, 4'hd, 4'hc, 4'h0, 4'hf, 4'h1, 4'h5, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h4, 4'h3, 4'h0, 4'hf, 4'h1, 4'h4, 4'h0 };
assign dw_0[893] = dw_0_893[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_894 = { 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h7, 4'h3, 4'h0, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h5, 4'h3, 4'hf, 4'h4, 4'h0, 4'hc, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h7, 4'h3, 4'h0, 4'hf, 4'h1, 4'h4, 4'h0 };
assign dw_0[894] = dw_0_894[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_895 = { 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h3, 4'h0, 4'h3, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h3, 4'h0, 4'h4, 4'h3, 4'hc, 4'h0, 4'h1, 4'hc, 4'h0, 4'hf, 4'h7, 4'h5, 4'h4, 4'h0, 4'h5, 4'h0, 4'hc, 4'hc, 4'hd, 4'hf, 4'h1, 4'h0, 4'hd, 4'h7, 4'h3, 4'h1, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'hd, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'h1, 4'h4, 4'h0 };
assign dw_0[895] = dw_0_895[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_896 = { 4'h3, 4'hd, 4'hc, 4'h1, 4'h0, 4'h3, 4'hf, 4'hd, 4'hc, 4'h1, 4'h1, 4'h0, 4'hc, 4'h3, 4'h3, 4'h1, 4'h3, 4'h3, 4'hd, 4'h3, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h0, 4'h4, 4'hd, 4'h7, 4'h0, 4'h3, 4'h1, 4'h0, 4'hf, 4'h3, 4'h4, 4'hc, 4'hc, 4'h1, 4'hc, 4'h1, 4'h0, 4'h3, 4'h4, 4'h5, 4'h4, 4'h0, 4'h4, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0 };
assign dw_0[896] = dw_0_896[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_897 = { 4'h3, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h1, 4'h5, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'hc, 4'hc, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h1, 4'h4, 4'h1, 4'h7, 4'h0, 4'h4, 4'h1, 4'h3, 4'hf, 4'h3, 4'h4, 4'hc, 4'h0, 4'hd, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'hc, 4'h1 };
assign dw_0[897] = dw_0_897[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_898 = { 4'hf, 4'hd, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'hd, 4'h1, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'hf, 4'h3, 4'hc, 4'hc, 4'h4, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'hf, 4'h1, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'hc, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h3, 4'h4, 4'hf, 4'hc, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h7, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0 };
assign dw_0[898] = dw_0_898[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_899 = { 4'hf, 4'hd, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hd, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'hc, 4'hf, 4'h3, 4'hc, 4'h4, 4'h3, 4'hd, 4'h0, 4'h0, 4'h1, 4'hd, 4'hf, 4'h1, 4'h0, 4'hc, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'hf, 4'h3, 4'h4, 4'hf, 4'h3, 4'hd, 4'h0, 4'h1, 4'h0, 4'h3, 4'h7, 4'h5, 4'h0, 4'hc, 4'h1, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0 };
assign dw_0[899] = dw_0_899[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_900 = { 4'hf, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'h1, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'hc, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'hf, 4'hc, 4'hd, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc };
assign dw_0[900] = dw_0_900[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_901 = { 4'hf, 4'hc, 4'hc, 4'h1, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'hd, 4'h1, 4'hc, 4'hc, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'hc, 4'h1, 4'h3, 4'hc, 4'hc, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'h5, 4'hc, 4'hf, 4'h0, 4'h3, 4'hd, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'hf, 4'h3, 4'h7, 4'hf, 4'hc, 4'hd, 4'h0, 4'hd, 4'h0, 4'h3, 4'h7, 4'h5, 4'h7, 4'h0, 4'h1, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0 };
assign dw_0[901] = dw_0_901[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_902 = { 4'hf, 4'hc, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'hd, 4'h1, 4'h0, 4'hc, 4'h3, 4'h3, 4'hd, 4'h0, 4'h1, 4'hd, 4'h0, 4'hf, 4'hc, 4'h0, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h5, 4'hc, 4'hf, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'hd, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h3, 4'hf, 4'hc, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h7, 4'h5, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0 };
assign dw_0[902] = dw_0_902[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_903 = { 4'hc, 4'hc, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'h4, 4'hc, 4'h1, 4'h3, 4'hc, 4'h0, 4'h3, 4'hd, 4'hd, 4'h1, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h4, 4'hc, 4'h4, 4'h7, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h3, 4'h4, 4'hc, 4'h0, 4'h1, 4'hc, 4'hd, 4'h0, 4'h3, 4'h7, 4'h5, 4'h4, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[903] = dw_0_903[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_904 = { 4'hf, 4'hd, 4'hc, 4'h1, 4'h0, 4'hc, 4'h3, 4'hf, 4'h5, 4'hd, 4'h1, 4'h3, 4'hf, 4'h0, 4'h3, 4'h1, 4'h1, 4'h1, 4'hd, 4'h1, 4'hc, 4'hf, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h3, 4'h4, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'hf, 4'h3, 4'h3, 4'hf, 4'hc, 4'h5, 4'h0, 4'hd, 4'h0, 4'h3, 4'h7, 4'h5, 4'h7, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[904] = dw_0_904[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_905 = { 4'hf, 4'hc, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h4, 4'hd, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'hd, 4'h1, 4'h0, 4'hd, 4'h1, 4'hf, 4'h0, 4'hc, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h5, 4'hc, 4'h4, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'hf, 4'hf, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc };
assign dw_0[905] = dw_0_905[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_906 = { 4'hf, 4'hd, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hd, 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h7, 4'hc, 4'h0, 4'h4, 4'h5, 4'hc, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h7, 4'hd, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'hc, 4'h5, 4'h0, 4'hc, 4'h0, 4'h3, 4'h7, 4'h5, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0 };
assign dw_0[906] = dw_0_906[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_907 = { 4'hf, 4'hf, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'h4, 4'hd, 4'h1, 4'h3, 4'hc, 4'h3, 4'h3, 4'h1, 4'h1, 4'h1, 4'hd, 4'h0, 4'hf, 4'hc, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'hd, 4'hf, 4'h0, 4'h4, 4'hc, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'hc, 4'h5, 4'h0, 4'hc, 4'h0, 4'h3, 4'h7, 4'h5, 4'h7, 4'hf, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc };
assign dw_0[907] = dw_0_907[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_908 = { 4'hf, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hd, 4'h3, 4'hf, 4'hc, 4'h0, 4'h3, 4'h1, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'hf, 4'h3, 4'h4, 4'hf, 4'hf, 4'h4, 4'hc, 4'hd, 4'h0, 4'h0, 4'h7, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0 };
assign dw_0[908] = dw_0_908[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_909 = { 4'hc, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hd, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'hc, 4'hc, 4'h4, 4'h7, 4'h1, 4'h0, 4'h0, 4'h5, 4'hc, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'h3, 4'hf, 4'h3, 4'h4, 4'hf, 4'hc, 4'h5, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3, 4'hc, 4'hc, 4'h4 };
assign dw_0[909] = dw_0_909[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_910 = { 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h7, 4'h3, 4'hc, 4'h3, 4'h0, 4'hd, 4'h0, 4'h3, 4'hf, 4'h3, 4'h3, 4'hc, 4'hf, 4'h4, 4'h4, 4'h1, 4'h0, 4'h4, 4'h5, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h3, 4'hf, 4'h3, 4'h4, 4'hf, 4'hc, 4'h4, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h3, 4'h5, 4'h0, 4'hf, 4'hc, 4'h0, 4'h5 };
assign dw_0[910] = dw_0_910[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_911 = { 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'hd, 4'h0, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h4, 4'h3, 4'hc, 4'h4, 4'hc, 4'h4, 4'hc, 4'h4, 4'h1, 4'h3, 4'hf, 4'h3, 4'h4, 4'hf, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h7, 4'h5, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0 };
assign dw_0[911] = dw_0_911[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_912 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'hc, 4'h4, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3, 4'h7, 4'h0, 4'h4, 4'h1, 4'h3, 4'h4, 4'h3, 4'h0, 4'h4, 4'h4, 4'hc, 4'h5, 4'h5, 4'h0, 4'hc, 4'h0, 4'hc, 4'hf, 4'h3, 4'hc, 4'h0, 4'hd, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h5, 4'h0, 4'hc, 4'h3, 4'hc, 4'h1 };
assign dw_0[912] = dw_0_912[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_913 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h7, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h4, 4'hc, 4'hc, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h5, 4'h3, 4'h3, 4'hc, 4'h4, 4'h1, 4'h3, 4'h4, 4'h7, 4'hc, 4'h4, 4'h5, 4'hc, 4'h5, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'hf, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1 };
assign dw_0[913] = dw_0_913[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_914 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'hc, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h5, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hd, 4'h1, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'hd, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0 };
assign dw_0[914] = dw_0_914[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_915 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h3, 4'h1, 4'h7, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'hc, 4'h4, 4'h7, 4'hc, 4'h0, 4'h0, 4'h4, 4'hf, 4'h3, 4'h1, 4'h4, 4'h4, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hd, 4'hc, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'hf, 4'h0, 4'hc, 4'hf };
assign dw_0[915] = dw_0_915[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_916 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h1, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h3, 4'h4, 4'h0, 4'h3, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'h1, 4'h0, 4'h4, 4'h1, 4'hf, 4'h4, 4'hc, 4'h0, 4'hd, 4'hc, 4'h5, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'h4, 4'hc, 4'h0, 4'h1, 4'hd, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3 };
assign dw_0[916] = dw_0_916[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_917 = { 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'hf, 4'h1, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'hd, 4'h3, 4'h3, 4'h3, 4'hf, 4'hc, 4'hc, 4'h4, 4'h4, 4'hf, 4'hc, 4'h0, 4'h0, 4'h7, 4'h3, 4'h3, 4'h1, 4'h4, 4'h4, 4'h1, 4'hf, 4'h4, 4'h0, 4'h1, 4'hd, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h5, 4'h1, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3 };
assign dw_0[917] = dw_0_917[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_918 = { 4'hc, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h1, 4'hf, 4'h3, 4'hc, 4'hf, 4'h4, 4'h1, 4'h3, 4'h0, 4'hf, 4'hf, 4'hc, 4'hc, 4'h4, 4'h4, 4'hc, 4'hc, 4'h0, 4'hc, 4'h7, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h4, 4'hc, 4'h0, 4'h5, 4'h3, 4'h4, 4'hc, 4'h0, 4'h1, 4'hf, 4'hc, 4'h0, 4'h0, 4'hd, 4'hc, 4'h3, 4'h4, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3 };
assign dw_0[918] = dw_0_918[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_919 = { 4'h3, 4'hc, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h1, 4'hf, 4'h0, 4'hc, 4'hf, 4'h4, 4'hd, 4'hd, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'hd, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h5, 4'hc, 4'h0, 4'h4, 4'h3, 4'h4, 4'hc, 4'h0, 4'h1, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hf, 4'h4, 4'h0, 4'h3, 4'h1, 4'h1, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3 };
assign dw_0[919] = dw_0_919[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_920 = { 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'h4, 4'h1, 4'h1, 4'h3, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'h1, 4'h3, 4'h1, 4'h1, 4'hf, 4'h0, 4'h0, 4'h5, 4'hc, 4'hc, 4'h5, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h7, 4'h0, 4'h3, 4'hd, 4'h1, 4'h0, 4'hf, 4'h3, 4'hc, 4'h3 };
assign dw_0[920] = dw_0_920[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_921 = { 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'hc, 4'h1, 4'h0, 4'hd, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'hd, 4'h1, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h4, 4'hf, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hd, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'h0, 4'h5, 4'hc, 4'h0, 4'h4, 4'h3, 4'h4, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'h5, 4'h0, 4'hd, 4'h0, 4'h3, 4'h7, 4'h0, 4'h0, 4'h1, 4'hd, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3 };
assign dw_0[921] = dw_0_921[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_922 = { 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h1, 4'hf, 4'h1, 4'hf, 4'hc, 4'hf, 4'hc, 4'h4, 4'hd, 4'h3, 4'h0, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h1, 4'hf, 4'h0, 4'h3, 4'h1, 4'hd, 4'h0, 4'h1, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h7, 4'h0, 4'h0, 4'h1, 4'hd, 4'h0, 4'hf, 4'hf, 4'hc, 4'hf };
assign dw_0[922] = dw_0_922[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_923 = { 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h4, 4'hc, 4'h0, 4'h1, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h3, 4'hd, 4'h0, 4'h4, 4'h1, 4'h3, 4'h5, 4'h0, 4'h4, 4'h0, 4'hc, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'h7, 4'h0, 4'hf, 4'h1, 4'hc, 4'h0, 4'hf, 4'hc, 4'hc, 4'hc };
assign dw_0[923] = dw_0_923[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_924 = { 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h7, 4'hc, 4'hf, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd, 4'h0, 4'h1, 4'h5, 4'h3, 4'h4, 4'h0, 4'h4, 4'h4, 4'hc, 4'h5, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'hf, 4'hc, 4'h0, 4'h4, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'hd, 4'h0, 4'hf, 4'hf, 4'hc, 4'hc };
assign dw_0[924] = dw_0_924[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_925 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'hc, 4'h0, 4'h7, 4'hf, 4'hf, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'hc, 4'h4, 4'h4, 4'hc, 4'h4, 4'h0, 4'h4, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'hc, 4'h5, 4'h1, 4'h1, 4'h3, 4'h3, 4'h0, 4'hf, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'hc, 4'h1, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0 };
assign dw_0[925] = dw_0_925[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_926 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'hf, 4'h3, 4'h1, 4'hc, 4'hc, 4'hc, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h7, 4'h5, 4'hc, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'hf, 4'h1, 4'h0, 4'hf, 4'h3, 4'h0, 4'h1 };
assign dw_0[926] = dw_0_926[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_927 = { 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h7, 4'hc, 4'h0, 4'hc, 4'h4, 4'h5, 4'h0, 4'h0, 4'hf, 4'h3, 4'h1, 4'hc, 4'h0, 4'hc, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h4, 4'h1, 4'h3, 4'h7, 4'h3, 4'h0, 4'h4, 4'h4, 4'hc, 4'h5, 4'h5, 4'h0, 4'hc, 4'h3, 4'hc, 4'hc, 4'hc, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h5, 4'h0, 4'hc, 4'hf, 4'h0, 4'h1 };
assign dw_0[927] = dw_0_927[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_928 = { 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'hf, 4'h5, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h4, 4'hf, 4'h1, 4'h1, 4'h1, 4'h1, 4'h4, 4'h7, 4'h1, 4'hc, 4'h5, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'h4, 4'hd, 4'h5, 4'h1, 4'h4, 4'h5, 4'h1, 4'h0, 4'h4, 4'h1, 4'h4, 4'h7, 4'h7, 4'h3, 4'hc, 4'h3, 4'h0, 4'h5, 4'hd, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h1, 4'h7, 4'h4, 4'h1 };
assign dw_0[928] = dw_0_928[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_929 = { 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'hd, 4'hd, 4'h1, 4'h0, 4'h4, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h7, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'hc, 4'h4, 4'hf, 4'h3, 4'h1, 4'h5, 4'h0, 4'h7, 4'h4, 4'h0, 4'h3, 4'h0, 4'h7, 4'h3, 4'h0, 4'hc, 4'h3, 4'h3, 4'h3, 4'hc, 4'hf, 4'h4, 4'h0, 4'hc, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h5, 4'h3, 4'h0, 4'h1 };
assign dw_0[929] = dw_0_929[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_930 = { 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1, 4'h1, 4'hd, 4'h0, 4'h4, 4'h0, 4'h7, 4'hc, 4'hc, 4'h3, 4'h1, 4'h0, 4'h7, 4'h7, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hd, 4'h3, 4'h1, 4'h3, 4'hc, 4'h3, 4'h0, 4'h5, 4'h4, 4'h7, 4'h7, 4'h0, 4'h3, 4'h0, 4'h7, 4'h4, 4'h1, 4'h0, 4'h7, 4'h4, 4'h3, 4'h3, 4'hf, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h5, 4'h0, 4'h4, 4'h1 };
assign dw_0[930] = dw_0_930[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_931 = { 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'hc, 4'hd, 4'h4, 4'h0, 4'hc, 4'h7, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'h1, 4'h4, 4'hf, 4'h0, 4'h0, 4'h4, 4'h7, 4'h4, 4'h7, 4'h0, 4'h3, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'h7, 4'h4, 4'h7, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1 };
assign dw_0[931] = dw_0_931[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_932 = { 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h3, 4'h3, 4'h7, 4'h7, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h7, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h4, 4'h7, 4'h4, 4'h3, 4'h3, 4'h7, 4'h4, 4'h0, 4'hd, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'hc, 4'hc, 4'h1, 4'h7, 4'h0, 4'h4, 4'h3, 4'h4, 4'h3 };
assign dw_0[932] = dw_0_932[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_933 = { 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'hd, 4'hc, 4'hd, 4'h5, 4'h4, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h3, 4'h3, 4'h4, 4'h0, 4'hc, 4'h0, 4'h3, 4'h4, 4'h0, 4'hc, 4'h1, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h5, 4'h7, 4'h4, 4'hf, 4'h7, 4'h7, 4'h4, 4'h1, 4'hd, 4'h4, 4'h4, 4'h3, 4'h3, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0 };
assign dw_0[933] = dw_0_933[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_934 = { 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h4, 4'h4, 4'h0, 4'h4, 4'h7, 4'hc, 4'h0, 4'h1, 4'h0, 4'h7, 4'h7, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h1, 4'h4, 4'hd, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h3, 4'h4, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h4, 4'h7, 4'h3, 4'h3, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h1, 4'h7, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0 };
assign dw_0[934] = dw_0_934[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_935 = { 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'hc, 4'hd, 4'h4, 4'h0, 4'hc, 4'h4, 4'h3, 4'hc, 4'h0, 4'h1, 4'hc, 4'h7, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hd, 4'hc, 4'h1, 4'h4, 4'hf, 4'h0, 4'h1, 4'h4, 4'h7, 4'h4, 4'h3, 4'h4, 4'hc, 4'h0, 4'h7, 4'h4, 4'h1, 4'h0, 4'h7, 4'h7, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h7, 4'h0, 4'h5, 4'h4, 4'h4, 4'hf };
assign dw_0[935] = dw_0_935[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_936 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'hd, 4'hc, 4'hd, 4'h7, 4'h0, 4'hc, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h4, 4'hd, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hd, 4'hf, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h4, 4'h4, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h7, 4'h7, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h1, 4'h7, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0 };
assign dw_0[936] = dw_0_936[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_937 = { 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'hd, 4'h3, 4'hc, 4'h0, 4'h7, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h7, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'hf, 4'h1, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h4, 4'hc, 4'h4, 4'h3, 4'h4, 4'h1, 4'hc, 4'h7, 4'h7, 4'h7, 4'h0, 4'hf, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'h1, 4'h7, 4'h0, 4'h5, 4'h4, 4'h4, 4'hf };
assign dw_0[937] = dw_0_937[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_938 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'hc, 4'hc, 4'h4, 4'h7, 4'h0, 4'h4, 4'h7, 4'h0, 4'h0, 4'h4, 4'h3, 4'h7, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'hd, 4'hc, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'hc, 4'h7, 4'h7, 4'h3, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h5, 4'h4, 4'h4, 4'h3 };
assign dw_0[938] = dw_0_938[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_939 = { 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'hd, 4'h0, 4'h7, 4'hc, 4'h7, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'hd, 4'hf, 4'h1, 4'h4, 4'hc, 4'h3, 4'h0, 4'h4, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'h3, 4'h7, 4'h7, 4'h7, 4'hc, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h3 };
assign dw_0[939] = dw_0_939[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_940 = { 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h7, 4'hc, 4'h7, 4'h3, 4'hc, 4'h0, 4'hd, 4'hc, 4'h7, 4'h7, 4'hd, 4'h4, 4'h7, 4'h3, 4'h1, 4'h0, 4'hd, 4'h1, 4'hc, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h4, 4'h4, 4'h4, 4'hd, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'h7, 4'h7, 4'h7, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'hf };
assign dw_0[940] = dw_0_940[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_941 = { 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h7, 4'h4, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'hc, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'hc, 4'h0, 4'hf, 4'h1, 4'h7, 4'hc, 4'h3, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'h4, 4'h7, 4'h7, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc, 4'h3, 4'hc, 4'hc, 4'h0, 4'h1, 4'h4, 4'h4, 4'h3 };
assign dw_0[941] = dw_0_941[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_942 = { 4'hc, 4'h7, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'hd, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h7, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h4, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'h0, 4'h1, 4'hf, 4'hc, 4'h1, 4'h4, 4'hc, 4'h3, 4'h1, 4'h7, 4'h0, 4'h7, 4'h4, 4'h4, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'hc, 4'hc, 4'hf, 4'hc, 4'hd, 4'h0, 4'h5, 4'h4, 4'h4, 4'hf };
assign dw_0[942] = dw_0_942[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_943 = { 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'hd, 4'hc, 4'h5, 4'h0, 4'h7, 4'h1, 4'h7, 4'hf, 4'h0, 4'h1, 4'h1, 4'hf, 4'h4, 4'h4, 4'hd, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'h5, 4'h7, 4'hc, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h7, 4'h7, 4'h3, 4'hc, 4'h7, 4'h0, 4'h1, 4'hd, 4'h3, 4'h0, 4'hc, 4'hd, 4'h0, 4'h1, 4'h5, 4'h4, 4'h3 };
assign dw_0[943] = dw_0_943[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_944 = { 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h4, 4'h3, 4'h4, 4'h5, 4'h4, 4'hc, 4'h0, 4'hc, 4'h7, 4'h0, 4'h7, 4'h0, 4'h1, 4'h3, 4'h7, 4'h0, 4'hd, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h4 };
assign dw_0[944] = dw_0_944[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_945 = { 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h4, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h5, 4'h7, 4'h4, 4'h5, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h7, 4'h0, 4'h1, 4'h3, 4'h3, 4'hd, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0 };
assign dw_0[945] = dw_0_945[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_946 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h4, 4'h1, 4'h0, 4'h1, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'hc, 4'h7, 4'h1, 4'h3, 4'h1, 4'h5, 4'h0, 4'h3, 4'hd, 4'h1, 4'hf, 4'h3, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h4, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h4, 4'h3, 4'h0, 4'h3, 4'hd, 4'hc, 4'h1 };
assign dw_0[946] = dw_0_946[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_947 = { 4'h4, 4'h7, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'h0, 4'h0, 4'hc, 4'h5, 4'h5, 4'h1, 4'h1, 4'h4, 4'h0, 4'h3, 4'h3, 4'h5, 4'h0, 4'h4, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h3, 4'h0, 4'h5, 4'h0, 4'h3, 4'h1, 4'h1, 4'hf, 4'hd, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h4, 4'h7, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0 };
assign dw_0[947] = dw_0_947[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_948 = { 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h5, 4'hc, 4'h1, 4'h5, 4'hc, 4'h0, 4'h5, 4'h0, 4'h5, 4'h3, 4'h0, 4'h3, 4'hc, 4'h5, 4'h0, 4'h5, 4'h3, 4'h0, 4'h5, 4'h4, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h3, 4'hc, 4'h5, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h1, 4'h0, 4'h4, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1 };
assign dw_0[948] = dw_0_948[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_949 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h3, 4'h1, 4'h4, 4'hc, 4'h0, 4'h5, 4'h1, 4'h5, 4'h7, 4'h0, 4'h3, 4'hd, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'hc, 4'h4, 4'h1, 4'h7, 4'h4, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h3, 4'h1, 4'h1, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h7, 4'h0, 4'h0, 4'h1, 4'hc, 4'h1 };
assign dw_0[949] = dw_0_949[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_950 = { 4'h4, 4'h4, 4'hc, 4'h1, 4'h0, 4'h4, 4'h5, 4'h3, 4'h1, 4'h5, 4'h3, 4'h4, 4'h5, 4'h5, 4'h1, 4'h7, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h4, 4'h7, 4'h4, 4'h5, 4'h0, 4'h3, 4'h1, 4'h1, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'h1, 4'h3, 4'h1, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'h5, 4'h4, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0 };
assign dw_0[950] = dw_0_950[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_951 = { 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h5, 4'hc, 4'h4, 4'h5, 4'h0, 4'h5, 4'h7, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h5, 4'h4, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'hc, 4'h7, 4'h4, 4'h7, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h4, 4'h1, 4'h0, 4'h5, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h3, 4'h0, 4'h4, 4'h1, 4'hc, 4'h5 };
assign dw_0[951] = dw_0_951[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_952 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'hc, 4'hd, 4'h4, 4'h3, 4'h4, 4'h5, 4'h0, 4'h1, 4'h7, 4'h4, 4'h3, 4'hc, 4'h5, 4'h0, 4'h4, 4'h7, 4'h0, 4'h5, 4'h4, 4'hc, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'hc, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'hd, 4'h0, 4'h1, 4'h1, 4'h4, 4'h4, 4'h1, 4'h1, 4'h4, 4'h4, 4'h0, 4'hc, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1 };
assign dw_0[952] = dw_0_952[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_953 = { 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'hd, 4'h1, 4'hf, 4'h0, 4'h5, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h7, 4'h4, 4'h5, 4'h5, 4'hc, 4'h0, 4'hc, 4'h0, 4'h4, 4'h7, 4'h0, 4'h5, 4'h0, 4'h7, 4'hd, 4'h1, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h5, 4'h1, 4'h0, 4'h5, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1 };
assign dw_0[953] = dw_0_953[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_954 = { 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'h0, 4'h1, 4'h7, 4'h1, 4'h0, 4'hc, 4'h5, 4'h4, 4'h5, 4'h7, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'hc, 4'h0, 4'h5, 4'h7, 4'h0, 4'h5, 4'h0, 4'h3, 4'hd, 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'h5, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h0 };
assign dw_0[954] = dw_0_954[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_955 = { 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h0, 4'h1, 4'h7, 4'h0, 4'h3, 4'hc, 4'h1, 4'h5, 4'h4, 4'h4, 4'h4, 4'h5, 4'h4, 4'hc, 4'h0, 4'hc, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h5, 4'h1, 4'hd, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'h0 };
assign dw_0[955] = dw_0_955[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_956 = { 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h3, 4'h0, 4'h1, 4'hc, 4'h4, 4'h5, 4'h0, 4'h5, 4'h7, 4'h0, 4'h0, 4'hd, 4'h1, 4'h1, 4'h4, 4'h7, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'h1, 4'h1, 4'h0, 4'h3, 4'h1, 4'h1, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'h0, 4'h4, 4'h1, 4'h1, 4'h5, 4'h1, 4'h0, 4'h1, 4'h3, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h4 };
assign dw_0[956] = dw_0_956[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_957 = { 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'h4, 4'h5, 4'hc, 4'h4, 4'h5, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0, 4'hc, 4'h4, 4'h5, 4'h4, 4'h7, 4'h4, 4'h5, 4'h5, 4'hc, 4'h0, 4'hf, 4'h3, 4'h4, 4'h3, 4'h4, 4'h4, 4'h0, 4'h3, 4'hd, 4'h1, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h7, 4'h1, 4'hc, 4'h5, 4'h1, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h4 };
assign dw_0[957] = dw_0_957[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_958 = { 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'h4, 4'h5, 4'h0, 4'h4, 4'h5, 4'h0, 4'h5, 4'h7, 4'h0, 4'h3, 4'h0, 4'h1, 4'h5, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'hc, 4'h3, 4'h4, 4'h3, 4'h5, 4'h4, 4'h0, 4'h0, 4'hd, 4'h1, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h7, 4'h1, 4'h3, 4'h5, 4'h1, 4'h1, 4'h1, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'h0 };
assign dw_0[958] = dw_0_958[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_959 = { 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'hf, 4'h0, 4'h3, 4'h0, 4'h1, 4'h5, 4'h5, 4'h0, 4'h4, 4'h5, 4'h0, 4'hc, 4'h0, 4'hf, 4'h7, 4'h5, 4'h3, 4'h0, 4'h5, 4'h3, 4'h3, 4'hd, 4'hd, 4'hf, 4'hd, 4'hc, 4'h1, 4'hc, 4'h3, 4'h7, 4'h1, 4'hc, 4'h4, 4'h5, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'hc, 4'h7, 4'hf, 4'h0, 4'h3, 4'h1, 4'hc, 4'h0 };
assign dw_0[959] = dw_0_959[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_960 = { 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'hf, 4'h1, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'hc, 4'h1, 4'h1, 4'h1, 4'hc, 4'h1, 4'hf, 4'h0, 4'hf, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'hd, 4'hf, 4'hc, 4'h1, 4'h0, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'hf, 4'h0, 4'h7, 4'h3, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'hd, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'hd };
assign dw_0[960] = dw_0_960[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_961 = { 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'hd, 4'h0, 4'hc, 4'h3, 4'h1, 4'h3, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'hc, 4'h0, 4'hf, 4'h3, 4'h3, 4'hc, 4'h7, 4'hd, 4'hc, 4'hd, 4'h3, 4'hf, 4'h0, 4'h1, 4'h5, 4'hc, 4'h4, 4'h7, 4'hc, 4'hf, 4'h1, 4'h4, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'hd };
assign dw_0[961] = dw_0_961[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_962 = { 4'h3, 4'hd, 4'h4, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'hc, 4'h1, 4'h3, 4'h0, 4'hd, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'hd, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h1, 4'h5, 4'hc, 4'h4, 4'h4, 4'hc, 4'h3, 4'h1, 4'h3, 4'h3, 4'h0, 4'h3, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1 };
assign dw_0[962] = dw_0_962[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_963 = { 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'hc, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'hf, 4'h1, 4'h0, 4'h1, 4'hd, 4'h0, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h3, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1 };
assign dw_0[963] = dw_0_963[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_964 = { 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'h1, 4'h0, 4'h1, 4'hc, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h4, 4'hd, 4'h0, 4'h1, 4'hf, 4'h0, 4'h3, 4'h4, 4'h5, 4'hf, 4'hc, 4'h4, 4'hc, 4'hf, 4'h1, 4'h4, 4'hf, 4'h0, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd };
assign dw_0[964] = dw_0_964[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_965 = { 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'h1, 4'h3, 4'h4, 4'h3, 4'hc, 4'h3, 4'hf, 4'h1, 4'h0, 4'h1, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h7, 4'hd, 4'h3, 4'h1, 4'h3, 4'h1, 4'hf, 4'h7, 4'h5, 4'hc, 4'h4, 4'h7, 4'hc, 4'h0, 4'hd, 4'h4, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h5, 4'h4, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1 };
assign dw_0[965] = dw_0_965[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_966 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'hc, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0, 4'hc, 4'h1, 4'hc, 4'h1, 4'hd, 4'h0, 4'h3, 4'h3, 4'hf, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h3, 4'h3, 4'h4, 4'h0, 4'hf, 4'hc, 4'h4, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'hf, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1 };
assign dw_0[966] = dw_0_966[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_967 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'h3, 4'hc, 4'hf, 4'hc, 4'h1, 4'h0, 4'h1, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'hd, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'hf, 4'h3, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1 };
assign dw_0[967] = dw_0_967[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_968 = { 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'h3, 4'h1, 4'h3, 4'hc, 4'h3, 4'hf, 4'h1, 4'h0, 4'h1, 4'hd, 4'h1, 4'h7, 4'h0, 4'hf, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'hc, 4'h1, 4'hf, 4'hc, 4'hf, 4'h0, 4'h4, 4'hf, 4'h3, 4'h5, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'hf, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h4, 4'h7, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1 };
assign dw_0[968] = dw_0_968[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_969 = { 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'h1, 4'h0, 4'h1, 4'hc, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h3, 4'h1, 4'hc, 4'h0, 4'h3, 4'h4, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hd };
assign dw_0[969] = dw_0_969[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_970 = { 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'h1, 4'hc, 4'h0, 4'h7, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h1, 4'hf, 4'h3, 4'h3, 4'h3, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hf, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h1 };
assign dw_0[970] = dw_0_970[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_971 = { 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'hc, 4'hc, 4'h0, 4'h3, 4'hc, 4'h3, 4'hc, 4'h1, 4'h0, 4'h1, 4'hd, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'hd, 4'h3, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hd, 4'h4, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'hc, 4'hd, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1 };
assign dw_0[971] = dw_0_971[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_972 = { 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'hf, 4'hc, 4'h1, 4'hf, 4'h0, 4'hc, 4'h0, 4'hf, 4'h1, 4'h0, 4'h1, 4'hd, 4'h1, 4'h3, 4'h0, 4'h3, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h7, 4'h0, 4'hf, 4'h0, 4'h4, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1 };
assign dw_0[972] = dw_0_972[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_973 = { 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'hf, 4'hc, 4'hd, 4'hf, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h3, 4'h1, 4'hc, 4'hf, 4'h1, 4'h1, 4'h5, 4'hf, 4'h0, 4'h7, 4'h0, 4'hf, 4'h1, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'h4, 4'h3, 4'hd, 4'h0, 4'hc, 4'h3, 4'h4, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0 };
assign dw_0[973] = dw_0_973[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_974 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h3, 4'hf, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h3, 4'h4, 4'hc, 4'h0, 4'h4, 4'hc, 4'h4, 4'hd, 4'h0, 4'hd, 4'hc, 4'h3, 4'h3, 4'h0, 4'h4, 4'hc, 4'h3, 4'h7, 4'hc, 4'hf, 4'h1, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'hd, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1 };
assign dw_0[974] = dw_0_974[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_975 = { 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'hd, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'hf, 4'h1, 4'h1, 4'h1, 4'hd, 4'h1, 4'hf, 4'h0, 4'h3, 4'h4, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'h4, 4'hc, 4'h4, 4'h3, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h7, 4'hf, 4'hc, 4'h4, 4'hc, 4'h1, 4'h0, 4'h0, 4'h7, 4'h5, 4'h4, 4'hd, 4'hc, 4'h0, 4'h3, 4'h4, 4'hc, 4'h3 };
assign dw_0[975] = dw_0_975[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_976 = { 4'h1, 4'h3, 4'h4, 4'h1, 4'h0, 4'h4, 4'h4, 4'h3, 4'h1, 4'h3, 4'h1, 4'h4, 4'hc, 4'h0, 4'h4, 4'hc, 4'hc, 4'h1, 4'hc, 4'h1, 4'h5, 4'h4, 4'h7, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h7, 4'h4, 4'h0, 4'h7, 4'h0, 4'h4, 4'h0, 4'h0, 4'h7, 4'h7, 4'h1, 4'hf, 4'h4, 4'h5, 4'h3, 4'h0, 4'hf, 4'h0, 4'h1, 4'hf, 4'hc, 4'hf, 4'h1, 4'hf, 4'h0, 4'h5, 4'h5, 4'hc, 4'h0 };
assign dw_0[976] = dw_0_976[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_977 = { 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'hc, 4'h4, 4'hd, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'hc, 4'h1, 4'hc, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h4, 4'h0, 4'h1, 4'hd, 4'h7, 4'hc, 4'h3, 4'h3, 4'h0, 4'h7, 4'h7, 4'h1, 4'h4, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'hf, 4'h0, 4'h1, 4'h7, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h5, 4'hc, 4'h3 };
assign dw_0[977] = dw_0_977[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_978 = { 4'h1, 4'h7, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'hf, 4'h1, 4'h0, 4'hd, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd, 4'h7, 4'h0, 4'h3, 4'h7, 4'h4, 4'h7, 4'h7, 4'h1, 4'h0, 4'h0, 4'h4, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'hc, 4'h0 };
assign dw_0[978] = dw_0_978[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_979 = { 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h5, 4'hd, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h5, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h1, 4'h3, 4'hc, 4'h3, 4'h3, 4'h4, 4'h4, 4'h7, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h4, 4'h4, 4'h0, 4'hf, 4'h0, 4'h4, 4'hf, 4'hd, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h3 };
assign dw_0[979] = dw_0_979[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_980 = { 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h3, 4'hc, 4'h4, 4'hc, 4'h4, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hc, 4'h0, 4'h5, 4'hc, 4'hd, 4'h0, 4'h7, 4'h3, 4'h4, 4'hf, 4'h1, 4'h4, 4'h3, 4'h5, 4'h0, 4'h0, 4'h4, 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'hd, 4'hf, 4'h3, 4'h0, 4'h0, 4'h5, 4'h1, 4'hc, 4'h0 };
assign dw_0[980] = dw_0_980[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_981 = { 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc, 4'h4, 4'h0, 4'h3, 4'h7, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h7, 4'hf, 4'h0, 4'hf, 4'h0, 4'h4, 4'h3, 4'h5, 4'h4, 4'hd, 4'h4, 4'h7, 4'h7, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0 };
assign dw_0[981] = dw_0_981[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_982 = { 4'h1, 4'h7, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h5, 4'hc, 4'h4, 4'h0, 4'hf, 4'h7, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h1, 4'hc, 4'h1, 4'h1, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h7, 4'h5, 4'h4, 4'h0, 4'h0, 4'h7, 4'h4, 4'h0, 4'hf, 4'h4, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0 };
assign dw_0[982] = dw_0_982[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_983 = { 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hd, 4'h1, 4'hd, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h1, 4'h1, 4'h7, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h7, 4'h5, 4'h0, 4'h0, 4'h1, 4'h3, 4'h4, 4'h1, 4'hf, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h1, 4'hf, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'h0 };
assign dw_0[983] = dw_0_983[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_984 = { 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h5, 4'hc, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'hf, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0, 4'h3, 4'h5, 4'h3, 4'h3, 4'h5, 4'h0, 4'h0, 4'h5, 4'h7, 4'h4, 4'h0, 4'hf, 4'h5, 4'h0, 4'h0, 4'h4, 4'hf, 4'h0, 4'h1, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[984] = dw_0_984[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_985 = { 4'h1, 4'h7, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h1, 4'h1, 4'hd, 4'h4, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h7, 4'hf, 4'h3, 4'h3, 4'h0, 4'h7, 4'h7, 4'h4, 4'h0, 4'h0, 4'h4, 4'h3, 4'h4, 4'h0, 4'hf, 4'h4, 4'h4, 4'h4, 4'h0, 4'hf, 4'h0, 4'h1, 4'h3, 4'hd, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h3 };
assign dw_0[985] = dw_0_985[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_986 = { 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h7, 4'h4, 4'h3, 4'h1, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hd, 4'h3, 4'h5, 4'h4, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3, 4'h5, 4'h0, 4'h0, 4'h4, 4'h3, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h5, 4'h3, 4'h1, 4'hf, 4'h0, 4'h3, 4'h0, 4'h5, 4'h1, 4'hc, 4'h0 };
assign dw_0[986] = dw_0_986[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_987 = { 4'h0, 4'h7, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'hf, 4'hd, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'h3, 4'h3, 4'h3, 4'h0, 4'h4, 4'h7, 4'h5, 4'h4, 4'h1, 4'h0, 4'h3, 4'h7, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'hc, 4'h3 };
assign dw_0[987] = dw_0_987[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_988 = { 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'hf, 4'h0, 4'h5, 4'hd, 4'h4, 4'h0, 4'h3, 4'h7, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h7, 4'h3, 4'h3, 4'h3, 4'h0, 4'h4, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'h4, 4'h4, 4'h4, 4'h4, 4'hf, 4'h0, 4'h1, 4'hf, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'hc, 4'h3 };
assign dw_0[988] = dw_0_988[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_989 = { 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'hf, 4'h0, 4'h1, 4'hd, 4'h1, 4'h4, 4'h3, 4'h4, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h5, 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h7, 4'h0, 4'h0, 4'h7, 4'h0, 4'h4, 4'h7, 4'h5, 4'h0, 4'h1, 4'h7, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h1, 4'hf, 4'hd, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0 };
assign dw_0[989] = dw_0_989[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_990 = { 4'h1, 4'h7, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'hf, 4'hc, 4'h5, 4'hd, 4'h4, 4'h1, 4'h3, 4'h7, 4'h4, 4'hf, 4'h1, 4'hd, 4'h1, 4'h5, 4'h4, 4'h0, 4'h4, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h7, 4'hd, 4'h3, 4'h3, 4'h0, 4'h4, 4'h7, 4'h1, 4'h0, 4'h1, 4'h7, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'h3 };
assign dw_0[990] = dw_0_990[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_991 = { 4'h1, 4'h7, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'hd, 4'h1, 4'hd, 4'h7, 4'h0, 4'h3, 4'h7, 4'hc, 4'hf, 4'h1, 4'hc, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h5, 4'h3, 4'h3, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h7, 4'h1, 4'h4, 4'hd, 4'h0, 4'h3, 4'h4, 4'h0, 4'hf, 4'h4, 4'h5, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'hf, 4'hd, 4'hc, 4'h4, 4'hc, 4'h0, 4'h4, 4'h5, 4'hc, 4'h0 };
assign dw_0[991] = dw_0_991[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_992 = { 4'h3, 4'hd, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'h1, 4'hd, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'hf, 4'h0, 4'hd, 4'h7, 4'hf, 4'h3, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'hf, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h7, 4'h5, 4'h7, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0 };
assign dw_0[992] = dw_0_992[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_993 = { 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h1, 4'h1, 4'h3, 4'hc, 4'hf, 4'h3, 4'h4, 4'hc, 4'h1, 4'hd, 4'h1, 4'hf, 4'h3, 4'hc, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h4, 4'hc, 4'hc, 4'h0, 4'h1, 4'hd, 4'h0, 4'h0, 4'h3, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0 };
assign dw_0[993] = dw_0_993[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_994 = { 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'h4, 4'hc, 4'h0, 4'hd, 4'h1, 4'hf, 4'hf, 4'h3, 4'h3, 4'h4, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'hf, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hf, 4'h0, 4'h4, 4'hd, 4'h3, 4'h4, 4'h0, 4'h4, 4'h3, 4'h4, 4'hc, 4'h3, 4'h5, 4'h3, 4'hf, 4'h3, 4'h7, 4'hc, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h5, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1 };
assign dw_0[994] = dw_0_994[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_995 = { 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'h4, 4'h3, 4'hf, 4'hc, 4'hd, 4'h0, 4'h3, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'hd, 4'h0, 4'hf, 4'hc, 4'h3, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h7, 4'hd, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'h0, 4'hf, 4'h5, 4'h0, 4'hf, 4'h3, 4'h4, 4'hf, 4'hf, 4'hc, 4'h0, 4'hd, 4'h0, 4'hc, 4'h3, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0 };
assign dw_0[995] = dw_0_995[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_996 = { 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h4, 4'h3, 4'h3, 4'h0, 4'hd, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'hf, 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'hf, 4'hf, 4'hc, 4'h3, 4'hd, 4'h3, 4'h7, 4'hc, 4'h7, 4'h0, 4'h5, 4'h0, 4'hc, 4'h5, 4'h3, 4'hf, 4'h3, 4'h7, 4'hc, 4'h0, 4'hc, 4'h1, 4'hd, 4'h0, 4'h0, 4'h3, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h1 };
assign dw_0[996] = dw_0_996[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_997 = { 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'hc, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h7, 4'hd, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h3, 4'h3, 4'hc, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h7, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc };
assign dw_0[997] = dw_0_997[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_998 = { 4'hf, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h1, 4'h3, 4'hc, 4'h3, 4'h3, 4'h5, 4'hf, 4'h0, 4'hc, 4'h1, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h7, 4'hf, 4'h3, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0 };
assign dw_0[998] = dw_0_998[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_999 = { 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h3, 4'hc, 4'h1, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'hc, 4'h1, 4'h1, 4'h3, 4'hf, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h3, 4'hd, 4'h3, 4'h4, 4'hc, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'h7, 4'h3, 4'h3, 4'h3, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h5, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[999] = dw_0_999[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1000 = { 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h3, 4'hc, 4'h1, 4'h3, 4'h3, 4'h3, 4'h3, 4'h1, 4'hd, 4'h1, 4'hd, 4'h1, 4'hf, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'hf, 4'hc, 4'h0, 4'h3, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h7, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h4, 4'hc, 4'h3, 4'h7, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[1000] = dw_0_1000[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1001 = { 4'hf, 4'hf, 4'hc, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'hc, 4'h1, 4'h0, 4'hf, 4'h3, 4'h3, 4'h4, 4'h0, 4'h1, 4'hd, 4'h1, 4'hf, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'h3, 4'h3, 4'h0, 4'hf, 4'h3, 4'h7, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h5, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[1001] = dw_0_1001[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1002 = { 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h3, 4'hd, 4'h1, 4'h3, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'hf, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h7, 4'hc, 4'h3, 4'h0, 4'hd, 4'h3, 4'h3, 4'h4, 4'hc, 4'h0, 4'h3, 4'h3, 4'hf, 4'h3, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0 };
assign dw_0[1002] = dw_0_1002[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1003 = { 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'h4, 4'hf, 4'h3, 4'hc, 4'h1, 4'h3, 4'h0, 4'h3, 4'h3, 4'h4, 4'hc, 4'h0, 4'hd, 4'h0, 4'hf, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h7, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h7, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0, 4'hc, 4'h4 };
assign dw_0[1003] = dw_0_1003[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1004 = { 4'h3, 4'hc, 4'hc, 4'h1, 4'h0, 4'hc, 4'h4, 4'h3, 4'hf, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'hd, 4'h1, 4'hf, 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'hf, 4'h0, 4'h7, 4'hc, 4'h3, 4'h7, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'hc, 4'hd, 4'h0, 4'h0, 4'h3, 4'h5, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0 };
assign dw_0[1004] = dw_0_1004[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1005 = { 4'h3, 4'hf, 4'hc, 4'h1, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h1, 4'hd, 4'h0, 4'h3, 4'h0, 4'hf, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'h5, 4'hc, 4'hf, 4'hc, 4'h4, 4'hc, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'hf, 4'h3, 4'h4, 4'hf, 4'hf, 4'h7, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0 };
assign dw_0[1005] = dw_0_1005[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1006 = { 4'h3, 4'hd, 4'hc, 4'h1, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3, 4'h3, 4'h3, 4'hf, 4'h5, 4'hf, 4'h0, 4'hd, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'hf, 4'h1, 4'h3, 4'hd, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h7, 4'hf, 4'hc, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0 };
assign dw_0[1006] = dw_0_1006[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1007 = { 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h4, 4'h3, 4'hf, 4'hc, 4'hd, 4'h3, 4'hc, 4'h3, 4'h3, 4'h5, 4'hf, 4'h0, 4'hd, 4'h0, 4'hf, 4'h0, 4'h3, 4'h4, 4'hd, 4'h0, 4'hc, 4'hc, 4'h1, 4'hf, 4'hc, 4'hc, 4'h3, 4'hc, 4'h0, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hf, 4'h3, 4'h7, 4'hf, 4'hc, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0 };
assign dw_0[1007] = dw_0_1007[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1008 = { 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'hf, 4'h1, 4'hf, 4'h4, 4'hc, 4'h0, 4'h3, 4'h4, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h5, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'h7, 4'h7, 4'hc, 4'h7, 4'h5, 4'hc, 4'h4, 4'hd, 4'h4, 4'h0, 4'h0, 4'h3, 4'h3, 4'h7, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h3, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1 };
assign dw_0[1008] = dw_0_1008[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1009 = { 4'hd, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'hc, 4'h3, 4'h3, 4'h3, 4'h4, 4'h7, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'hc, 4'h3, 4'h3, 4'h3, 4'h4, 4'hc, 4'h7, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h7, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1 };
assign dw_0[1009] = dw_0_1009[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1010 = { 4'hd, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h0, 4'h3, 4'hf, 4'h4, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h3, 4'hf, 4'h4, 4'hc, 4'h7, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1 };
assign dw_0[1010] = dw_0_1010[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1011 = { 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h4, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc, 4'h1, 4'h0, 4'hf, 4'hf, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1 };
assign dw_0[1011] = dw_0_1011[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1012 = { 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'hf, 4'h1, 4'hc, 4'h4, 4'h3, 4'hd, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h3, 4'h1, 4'hd, 4'h3, 4'h1, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'hd, 4'h4, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[1012] = dw_0_1012[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1013 = { 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'h0, 4'h3, 4'hf, 4'h4, 4'h7, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'hc, 4'h1, 4'h1, 4'h7, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hd, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1 };
assign dw_0[1013] = dw_0_1013[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1014 = { 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'hd, 4'hd, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'hd, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'hc, 4'h3, 4'h1, 4'hf, 4'h4, 4'h1, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'h0, 4'hc, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hf, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0 };
assign dw_0[1014] = dw_0_1014[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1015 = { 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'hf, 4'h4, 4'hc, 4'h0, 4'h3, 4'h1, 4'hc, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'hf, 4'h1, 4'hc, 4'h0, 4'h1, 4'hc, 4'h4, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h5, 4'h4, 4'h0, 4'h1, 4'h3, 4'h0, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'hf, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3 };
assign dw_0[1015] = dw_0_1015[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1016 = { 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'h0, 4'h4, 4'h1, 4'hc, 4'h1, 4'hc, 4'h3, 4'h1, 4'hf, 4'h4, 4'h5, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'h3, 4'h7, 4'h4, 4'h1, 4'hf, 4'h0, 4'h0, 4'h7, 4'hc, 4'hc, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[1016] = dw_0_1016[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1017 = { 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'hd, 4'h0, 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'h1, 4'hd, 4'h3, 4'h1, 4'hc, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h4, 4'h1, 4'hf, 4'h0, 4'h0, 4'h4, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[1017] = dw_0_1017[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1018 = { 4'hc, 4'h7, 4'h4, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h1, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0, 4'h3, 4'hc, 4'hd, 4'h1, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'hd, 4'hc, 4'h3, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hc, 4'h4, 4'h4, 4'h3, 4'hc, 4'h3, 4'h3, 4'h7, 4'h1, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[1018] = dw_0_1018[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1019 = { 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'h3, 4'hf, 4'h4, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'hc, 4'hd, 4'hc, 4'h0, 4'h1, 4'hc, 4'h4, 4'h0, 4'h4, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[1019] = dw_0_1019[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1020 = { 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'hf, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'hd, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'hf, 4'h1, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'h4, 4'h0, 4'h4, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0 };
assign dw_0[1020] = dw_0_1020[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1021 = { 4'hd, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'hd, 4'hc, 4'h4, 4'h0, 4'h3, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'h3, 4'hf, 4'h4, 4'h3, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'h4, 4'hc, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'hc, 4'h7, 4'h4, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'h3, 4'hf, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1 };
assign dw_0[1021] = dw_0_1021[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1022 = { 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'hd, 4'hc, 4'h0, 4'h1, 4'h3, 4'h4, 4'h1, 4'h3, 4'h0, 4'h3, 4'hd, 4'h0, 4'h0, 4'h3, 4'hc, 4'h5, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h3, 4'h4, 4'hc, 4'h7, 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'h3, 4'h3, 4'hd, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1 };
assign dw_0[1022] = dw_0_1022[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1023 = { 4'hc, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'hc, 4'h4, 4'h0, 4'h3, 4'h0, 4'h7, 4'hc, 4'h1, 4'h0, 4'hf, 4'h0, 4'h5, 4'h0, 4'hc, 4'hc, 4'h4, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'hc, 4'h1, 4'h1, 4'hc, 4'h3, 4'h0, 4'h7, 4'hc, 4'h7, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h3, 4'hd, 4'h0, 4'h3, 4'h4, 4'h4, 4'h1 };
assign dw_0[1023] = dw_0_1023[d0_cntr];
