localparam D0_IN_SIZE = 2;
localparam D0_BW_W = 2;
localparam D0_SHIFT = 0;
localparam LOG2_D0_CYC = 9;
localparam D0_CYC = 512;
localparam D0_CH = 128;
reg [LOG2_D0_CYC-1:0] d0_cntr;
wire [D0_CH-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0;
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_0 = { 4'h5, 4'h4, 4'h0, 4'h0, 4'hc, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'hd, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h1, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h3, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'h3, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h5, 4'h4, 4'h0, 4'h3, 4'hf, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h5, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h0, 4'h3, 4'h3, 4'hf, 4'h3, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'hc, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'hf, 4'h5, 4'h3, 4'h3, 4'h3, 4'hf, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'hf, 4'h3, 4'hf, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'h4, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf };
assign dw_0[0] = dw_0_0[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_1 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h1, 4'h0, 4'h4, 4'h1, 4'h4, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h1, 4'h0, 4'h5, 4'h0, 4'h4, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'h4, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h3, 4'hc, 4'hc, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h4, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h1, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h5, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0 };
assign dw_0[1] = dw_0_1[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_2 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[2] = dw_0_2[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_3 = { 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'hf, 4'h0, 4'hc, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'hc, 4'hc, 4'hf, 4'hf, 4'hc, 4'h5, 4'h4, 4'h4, 4'h5, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'hc, 4'hc, 4'hc, 4'h0, 4'h3, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h4, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h3, 4'hc, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h5, 4'h4, 4'h1, 4'h1, 4'h0, 4'h1, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h3, 4'hc, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h1, 4'hc, 4'hc, 4'hf, 4'h3, 4'hc, 4'h3, 4'hc, 4'h3, 4'h3, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'h1, 4'h5, 4'h0, 4'h5, 4'h0, 4'h4, 4'h3, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h5, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h4, 4'h1, 4'h1, 4'h0, 4'h4, 4'h3, 4'h1, 4'h5, 4'h4, 4'h1, 4'h0, 4'h4, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h3, 4'hc, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hc, 4'h3, 4'h3, 4'h3, 4'hf, 4'h0, 4'h1, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h4, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h5, 4'hd, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[3] = dw_0_3[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_4 = { 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h5, 4'h1, 4'h5, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h1, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h1, 4'h5, 4'h0, 4'h1, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h1, 4'h4, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h4, 4'h5, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'hf, 4'h0, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'hc, 4'h0, 4'h3, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf };
assign dw_0[4] = dw_0_4[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_5 = { 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h1, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'hc, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'hf, 4'hf, 4'hc, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h4, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h7, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1 };
assign dw_0[5] = dw_0_5[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_6 = { 4'hc, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'hf, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h4, 4'h1, 4'h5, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h4, 4'h5, 4'h1, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'h1, 4'h5, 4'h4, 4'h1, 4'h4, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'h0, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'h3, 4'h0, 4'h3, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h4, 4'h1, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h5, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'h4, 4'h3, 4'h3, 4'h0, 4'h1, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h1, 4'h5, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'h3, 4'h3, 4'hc, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'hf, 4'h3, 4'h1, 4'h3, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h3, 4'h3, 4'hc, 4'hf, 4'hf, 4'h4, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'h3, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h5, 4'h4, 4'h5, 4'h4, 4'h1, 4'h5 };
assign dw_0[6] = dw_0_6[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_7 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h0, 4'h4, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'hf, 4'hc, 4'h3, 4'hc, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h0, 4'h5, 4'h1, 4'h5, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h1, 4'h4, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h3, 4'hf, 4'h3, 4'hf, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h5, 4'h0, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[7] = dw_0_7[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_8 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[8] = dw_0_8[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_9 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[9] = dw_0_9[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_10 = { 4'h5, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h5, 4'h1, 4'h0, 4'h5, 4'h4, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h5, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h5, 4'h5, 4'h1, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0, 4'hf, 4'h4, 4'h1, 4'h4, 4'h1, 4'h5, 4'h4, 4'h5, 4'h1, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'hf, 4'h0, 4'h5, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'h4, 4'h0, 4'h1, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'hd, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h4, 4'h1, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h4, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'hf, 4'h3, 4'h4, 4'h5, 4'h0, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'hf, 4'hc, 4'h3, 4'hc, 4'hf, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'hd, 4'h1, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'hc, 4'h4, 4'h4, 4'h0, 4'h7, 4'h0, 4'h3, 4'h5, 4'h5, 4'h1, 4'h1, 4'hc, 4'h3, 4'h3, 4'h3, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'hc, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0 };
assign dw_0[10] = dw_0_10[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_11 = { 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'hf, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h4, 4'h3, 4'hf, 4'hc, 4'h0, 4'h3, 4'hf, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h1, 4'h1, 4'h1, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'h1, 4'h1, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0 };
assign dw_0[11] = dw_0_11[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_12 = { 4'hf, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h5, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h1, 4'h0, 4'h7, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h5, 4'h5, 4'h4, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'hf, 4'hf, 4'h0, 4'h1, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'h1, 4'h4, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h5, 4'h5, 4'h0, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h3, 4'h3, 4'h5, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h1, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h7, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1 };
assign dw_0[12] = dw_0_12[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_13 = { 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h1, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h5, 4'h3, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h4, 4'h1, 4'h5, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf };
assign dw_0[13] = dw_0_13[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_14 = { 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'hc, 4'h4, 4'h0, 4'h3, 4'h3, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'h3, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h0, 4'h3, 4'h3, 4'h4, 4'h3, 4'h0, 4'h3, 4'h3, 4'hf, 4'hc, 4'hf, 4'h3, 4'hc, 4'hf, 4'h3, 4'h3, 4'h3, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h5, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h1, 4'h1, 4'h3, 4'h1, 4'h5, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'h0, 4'h4, 4'h1, 4'h1, 4'h4, 4'hd, 4'h4, 4'h1, 4'h5, 4'h1, 4'h5, 4'h0, 4'h4, 4'h1, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h3, 4'h3, 4'h3, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h4, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h5, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h0, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'hc, 4'hd, 4'hd, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h0, 4'h5, 4'h4, 4'h4, 4'h5, 4'h0, 4'h5, 4'h1, 4'h4, 4'h1, 4'h4, 4'h4, 4'h1, 4'h0, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'hc, 4'hd, 4'h0, 4'h0 };
assign dw_0[14] = dw_0_14[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_15 = { 4'hc, 4'h0, 4'h3, 4'hf, 4'h0, 4'hc, 4'hf, 4'h3, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'hc, 4'h3, 4'h3, 4'hf, 4'h3, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5, 4'h4, 4'h4, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h4, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'hc, 4'h3, 4'h3, 4'h4, 4'h4, 4'h4, 4'h0, 4'h1, 4'h5, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h5, 4'h4, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h1, 4'h1, 4'h0, 4'h4, 4'h5, 4'h1, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'hc, 4'h3, 4'hc, 4'h0, 4'hc, 4'hc, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h4, 4'h3, 4'hc, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h5, 4'h1, 4'h1, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h5, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'h1, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h0, 4'hd, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'hf, 4'hf, 4'h3, 4'h3, 4'h3, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h0, 4'hd, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'hc, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'h3, 4'hf, 4'hc, 4'h4, 4'h5, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h1, 4'h0, 4'h5, 4'h0, 4'hc, 4'h4, 4'h0, 4'h1, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h3, 4'hf, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h0, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0 };
assign dw_0[15] = dw_0_15[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_16 = { 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'hf, 4'h3, 4'h1, 4'h0, 4'h1, 4'h5, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h3, 4'hc, 4'hf, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h5, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h5, 4'h3, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'hc, 4'h3, 4'hc, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'hc, 4'h1, 4'h5, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h4, 4'hf, 4'hc, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'h3, 4'h3, 4'h0, 4'hc, 4'hc, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'hf, 4'hc, 4'h3, 4'hc, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf };
assign dw_0[16] = dw_0_16[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_17 = { 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h1, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'hc, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'hf, 4'h3, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h0, 4'h4, 4'h1, 4'h5, 4'h1, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h5, 4'h5, 4'h0, 4'h4, 4'h5, 4'h5, 4'h4, 4'h4, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'hf, 4'hc, 4'hc, 4'hf, 4'hc, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'hf, 4'h0, 4'h5, 4'h4, 4'h0, 4'h4, 4'h1, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h5, 4'h1, 4'h4, 4'h4, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'h5, 4'h4, 4'h0, 4'h4, 4'hc, 4'h0, 4'hf, 4'h4, 4'hc, 4'h1, 4'h0, 4'hc, 4'h4, 4'h4, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h1, 4'hf, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'h7, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hc, 4'h0, 4'h3, 4'h3, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h7, 4'h5, 4'h5, 4'h0, 4'h4, 4'h5, 4'h4, 4'h1, 4'h1, 4'h5, 4'h1, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'hc, 4'h1, 4'h1, 4'h4, 4'h1, 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h3, 4'hf, 4'h3, 4'h0, 4'hc, 4'hf, 4'h0 };
assign dw_0[17] = dw_0_17[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_18 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h1, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h1, 4'h1, 4'h3, 4'h7, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h7, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'h3, 4'h3, 4'hf, 4'hc, 4'hf, 4'h4, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h0, 4'h5, 4'h5, 4'h1, 4'h0, 4'h4, 4'h5, 4'h1, 4'h1, 4'h0, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'hd, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h5, 4'h4, 4'h7, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'hf, 4'h3, 4'hc, 4'hf, 4'h3, 4'h3, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h4, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'hd, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'hd, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h4, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0 };
assign dw_0[18] = dw_0_18[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_19 = { 4'hf, 4'hf, 4'h1, 4'h5, 4'h5, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'hf, 4'h3, 4'h4, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'h4, 4'h1, 4'h5, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'hf, 4'h3, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'hf, 4'h3, 4'hc, 4'h3, 4'h3, 4'hf, 4'h3, 4'h5, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h5, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'hc, 4'h3, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h3, 4'h5, 4'h5, 4'h1, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h4, 4'h1, 4'hc, 4'h0, 4'h1, 4'h5, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'h4, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h4, 4'h1, 4'hc, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h4, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'hf, 4'h3, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0, 4'h5, 4'h0, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'hc, 4'hf, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h7, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd, 4'h1, 4'h1, 4'h1, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h5, 4'h1, 4'h1, 4'h1, 4'h1, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hc, 4'hc, 4'hc };
assign dw_0[19] = dw_0_19[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_20 = { 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'hf, 4'hf, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'h3, 4'hf, 4'h0, 4'hc, 4'hf, 4'hc, 4'hf, 4'h7, 4'hf, 4'hf, 4'h3, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'hf, 4'h3, 4'h3, 4'hf, 4'h3, 4'hc, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h0, 4'hc, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'h3, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'h3, 4'h3, 4'h3, 4'hf, 4'hc, 4'hc, 4'hc, 4'hc, 4'h3, 4'h3, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h1, 4'h5, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h5, 4'h4, 4'h0, 4'h4, 4'h5, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'h1, 4'h4, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[20] = dw_0_20[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_21 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[21] = dw_0_21[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_22 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[22] = dw_0_22[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_23 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h4, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h0, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[23] = dw_0_23[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_24 = { 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h5, 4'h0, 4'h1, 4'h1, 4'h1, 4'h5, 4'h4, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h4, 4'h0, 4'h1, 4'h1, 4'h1, 4'h4, 4'h1, 4'h3, 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h1, 4'h5, 4'h1, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h3, 4'h1, 4'h1, 4'h4, 4'h1, 4'h4, 4'h5, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hc, 4'hc, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h0, 4'h1, 4'h1, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h5, 4'h1, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'hc, 4'h0, 4'h4, 4'hf, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h4, 4'h4, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h1, 4'h1, 4'h5, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'hc, 4'h1, 4'hf, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'hd, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'hf, 4'h3, 4'hd, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h1, 4'h5, 4'h1, 4'h4, 4'h0, 4'h4, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'h1, 4'h4, 4'hc, 4'h4, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h7, 4'h3, 4'h7, 4'hc, 4'h3, 4'h3, 4'hd, 4'h1, 4'h5, 4'h0, 4'h4, 4'h5, 4'h4, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h3, 4'hf, 4'h3, 4'hc, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hc, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h4, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[24] = dw_0_24[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_25 = { 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h5, 4'h1, 4'h4, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'h3, 4'hf, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h4, 4'h4, 4'h4, 4'h0, 4'h5, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'h0, 4'h3, 4'hf, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h5, 4'h5, 4'h0, 4'h0, 4'h5, 4'h1, 4'h1, 4'h5, 4'h1, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'hf, 4'h3, 4'hc, 4'h3, 4'hf, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'hf, 4'hc, 4'h1, 4'h4, 4'h1, 4'h0, 4'h5, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'hf, 4'hc, 4'hd, 4'h1, 4'h3, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'hf, 4'hc, 4'hc, 4'hc, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h0, 4'h5, 4'h5, 4'h4, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'hd, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'hf, 4'hf, 4'h3, 4'h0, 4'h3, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'h5, 4'h4, 4'h4, 4'h5, 4'h1, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h4, 4'h1, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0 };
assign dw_0[25] = dw_0_25[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_26 = { 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h5, 4'h5, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'h4, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h5, 4'h1, 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h4, 4'h4, 4'h1, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'h1, 4'h4, 4'h1, 4'h1, 4'h4, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h0, 4'h5, 4'h4, 4'h0, 4'h5, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf };
assign dw_0[26] = dw_0_26[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_27 = { 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h5, 4'h4, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h3, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h5, 4'h4, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h4, 4'h1, 4'h5, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'h3, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'hc, 4'h4, 4'h4, 4'h3, 4'h0, 4'hf, 4'h0, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'h3, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h5, 4'h1, 4'h5, 4'h1, 4'h4, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'h3, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'h3, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf };
assign dw_0[27] = dw_0_27[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_28 = { 4'h0, 4'hc, 4'hf, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h0, 4'h4, 4'hc, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'h5, 4'h4, 4'h0, 4'h5, 4'h1, 4'h3, 4'h1, 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'h4, 4'h5, 4'h0, 4'h1, 4'h1, 4'h1, 4'h3, 4'h3, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'h1, 4'h1, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'hc, 4'hf, 4'h3, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'hc, 4'h3, 4'h3, 4'h3, 4'hc, 4'h3, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'h4, 4'h5, 4'h4, 4'h1, 4'h0, 4'h5, 4'h5, 4'h4, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'h1, 4'h5, 4'h5, 4'h4, 4'hc, 4'h0, 4'h1, 4'h4, 4'h1, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'h3, 4'h3, 4'h0, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'hf, 4'h5, 4'h5, 4'h0, 4'h1, 4'h5, 4'h4, 4'h0, 4'h4, 4'h3, 4'h3, 4'hf, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h1, 4'h7, 4'h1, 4'h5, 4'h1, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h3, 4'h3, 4'h3, 4'h4, 4'hf, 4'h5, 4'h5, 4'h4, 4'h0, 4'h3, 4'h5, 4'h0, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'hf, 4'h0, 4'h3, 4'h3, 4'hc, 4'h3, 4'hf, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h7, 4'hf, 4'h0, 4'hf, 4'hc, 4'hc, 4'hf, 4'hc, 4'h0, 4'h4, 4'h1, 4'h4, 4'h5, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'h7, 4'h3, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'h3, 4'h3, 4'hc, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h1, 4'h4, 4'h5, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hc, 4'hc, 4'h1, 4'h4, 4'h0, 4'hc, 4'h4, 4'h7, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4 };
assign dw_0[28] = dw_0_28[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_29 = { 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h4, 4'h4, 4'h1, 4'h0, 4'hf, 4'hf, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h0, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'hc, 4'hc, 4'h3, 4'hc, 4'h3, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h3, 4'hc, 4'hc, 4'h7, 4'hc, 4'h0, 4'h3, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h3, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h5, 4'h4, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'hf, 4'h1, 4'h3, 4'hf, 4'h0, 4'h4, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h0, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h1, 4'h4, 4'h5, 4'h0, 4'h5, 4'h5, 4'h0, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'hf, 4'h3, 4'h3, 4'h0, 4'h3, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h3, 4'hf, 4'hf, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'hf, 4'h3, 4'hf, 4'hc, 4'h4, 4'h0, 4'h3, 4'h1, 4'h5, 4'h4, 4'h4, 4'h5, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'hd, 4'h0, 4'hc, 4'h3, 4'h0, 4'hd, 4'hc, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'hf, 4'h3, 4'h0, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h7, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h4, 4'h5, 4'h4, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h4, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0 };
assign dw_0[29] = dw_0_29[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_30 = { 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'h3, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h0, 4'h4, 4'hf, 4'hc, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'h3, 4'hc, 4'hf, 4'hc, 4'h3, 4'hf, 4'h3, 4'h3, 4'h3, 4'hf, 4'h3, 4'hf, 4'hc, 4'h1, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'hc, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'hf, 4'hc, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'h0, 4'hc, 4'h0, 4'h1, 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'h1, 4'h4, 4'h4, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'hc, 4'hf };
assign dw_0[30] = dw_0_30[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_31 = { 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'h4, 4'h1, 4'h4, 4'h4, 4'h1, 4'h0, 4'h4, 4'h1, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'hf, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hf, 4'h3, 4'hc, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h3, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h5, 4'h1, 4'h4, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h4, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h1, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h3, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'hc, 4'hc, 4'h0, 4'hc, 4'hf, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0 };
assign dw_0[31] = dw_0_31[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_32 = { 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'hc, 4'h3, 4'hf, 4'h1, 4'h4, 4'h4, 4'h4, 4'h4, 4'h0, 4'h4, 4'h5, 4'hc, 4'h3, 4'hf, 4'hc, 4'hc, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h1, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'h0, 4'hf, 4'hc, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'hf, 4'h1, 4'h4, 4'h1, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'hf, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'h1, 4'h5, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h5, 4'h1, 4'h0, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h1, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'hc, 4'hf, 4'h0, 4'hf, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h5, 4'h0, 4'hc, 4'h3, 4'hf, 4'h3, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf };
assign dw_0[32] = dw_0_32[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_33 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'h3, 4'h3, 4'h3, 4'hf, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h7, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'hc, 4'hf, 4'hc, 4'hf, 4'h3, 4'hc, 4'h0, 4'hc, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h1, 4'h0, 4'h1, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hc, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hc, 4'hc, 4'hc, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h4, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'hf, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h1, 4'h5, 4'h4, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h7, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0 };
assign dw_0[33] = dw_0_33[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_34 = { 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'hf, 4'hc, 4'h3, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h1, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'hf, 4'h1, 4'hc, 4'h3, 4'h3, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'h0, 4'h3, 4'h4, 4'hc, 4'h0, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h1, 4'h5, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h5, 4'h4, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'h4, 4'h4, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'hd, 4'h4, 4'h0, 4'h5, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'hf, 4'h3, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'hc, 4'h3, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'h3, 4'hc, 4'h3, 4'hf, 4'h3, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'hc, 4'hc, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'h3, 4'hc, 4'hc, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'h5, 4'hc, 4'h1, 4'h1, 4'h5, 4'h5, 4'h3, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'h1, 4'h1, 4'h4, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h0 };
assign dw_0[34] = dw_0_34[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_35 = { 4'h0, 4'hf, 4'h3, 4'hc, 4'h3, 4'h1, 4'h3, 4'hc, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'h4, 4'h0, 4'h3, 4'h1, 4'h1, 4'h1, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'hd, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h5, 4'h5, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h1, 4'h5, 4'h0, 4'h4, 4'hd, 4'h5, 4'h4, 4'h5, 4'hf, 4'h1, 4'h4, 4'h0, 4'hf, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'hf, 4'hf, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h1, 4'h1, 4'h1, 4'h1, 4'h0, 4'h5, 4'hd, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'hf, 4'hf, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'h3, 4'hd, 4'hc, 4'h0, 4'h4, 4'h1, 4'hf, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'hf, 4'hc, 4'hc, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h4, 4'h4, 4'h0, 4'h5, 4'h0, 4'h4, 4'h5, 4'h1, 4'hf, 4'h3, 4'hf, 4'hc, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'hd, 4'h3, 4'h1, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h1, 4'hf, 4'h0, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h3, 4'h4, 4'hc, 4'hd, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h5, 4'h4, 4'h5, 4'h1, 4'h1, 4'h5, 4'h3, 4'hc, 4'h3, 4'h0, 4'hc, 4'hf, 4'hf, 4'h3, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'h4, 4'h1, 4'h5, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h4, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'hf, 4'h3, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h1, 4'h4, 4'h5, 4'h4, 4'h5, 4'h4, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h3, 4'h5, 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'h5, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h3, 4'hc, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'h4, 4'h4, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'hc, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5 };
assign dw_0[35] = dw_0_35[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_36 = { 4'h3, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h1, 4'h1, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'hf, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'hf, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[36] = dw_0_36[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_37 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[37] = dw_0_37[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_38 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h1, 4'h5, 4'h0, 4'h5, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'hc, 4'h3, 4'hc, 4'h3, 4'h1, 4'h0, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hd, 4'h4, 4'h4, 4'h1, 4'h4, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h1, 4'h4, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'h1, 4'h4, 4'h1, 4'h4, 4'h4, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h5, 4'h5, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h4, 4'h1, 4'h5, 4'h1, 4'h5, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'h7, 4'h0, 4'h5, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hd, 4'h5, 4'h1, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'hc, 4'hc, 4'hf, 4'h3, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'hc, 4'hd, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5 };
assign dw_0[38] = dw_0_38[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_39 = { 4'h0, 4'h4, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'hf, 4'hc, 4'h0, 4'hf, 4'hc, 4'hf, 4'h5, 4'h5, 4'h4, 4'h4, 4'h4, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h1, 4'h1, 4'hc, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'hc, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h5, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'h1, 4'h0, 4'h5, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h1, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'hf, 4'h4, 4'h0, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'h3, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h1, 4'h4, 4'h0, 4'h5, 4'h1, 4'h0, 4'h1, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h1, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'h3, 4'hf, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h4, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'hd, 4'h3, 4'hc, 4'hf, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h5, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h3, 4'hf, 4'hf, 4'h0, 4'h3, 4'hf, 4'hf, 4'hc, 4'h3, 4'hc, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'hc, 4'hc, 4'h3, 4'h4, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h5, 4'h1, 4'h4, 4'h1, 4'h1, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'hc, 4'hc, 4'hf, 4'h0, 4'hc, 4'hf, 4'h0 };
assign dw_0[39] = dw_0_39[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_40 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'h1, 4'h1, 4'h4, 4'h4, 4'h3, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h1, 4'hf, 4'hc, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h4, 4'h7, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h5, 4'h4, 4'h0, 4'h5, 4'h0, 4'h1, 4'h5, 4'hc, 4'h0, 4'h4, 4'h1, 4'h5, 4'h5, 4'h1, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h3, 4'hf, 4'hc, 4'hc, 4'hc, 4'h7, 4'h0, 4'hc, 4'h3, 4'hc, 4'h3, 4'h3, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'hc, 4'h0, 4'hc, 4'hf, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'h4, 4'h5, 4'h4, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'hc, 4'h3, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'hc, 4'h1, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'h1, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'hf, 4'h3, 4'hf, 4'hc, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'hf, 4'h0, 4'hc, 4'hf, 4'hc, 4'h0, 4'h3, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'h4, 4'h1, 4'h5, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h3, 4'h0, 4'h1, 4'h7, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3 };
assign dw_0[40] = dw_0_40[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_41 = { 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'hc, 4'h3, 4'h3, 4'h3, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'hf, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'h3, 4'h1, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h5, 4'h1, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h5, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'hf, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h5, 4'h5 };
assign dw_0[41] = dw_0_41[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_42 = { 4'h5, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'h1, 4'h5, 4'h4, 4'h0, 4'hf, 4'hc, 4'hc, 4'h1, 4'h5, 4'h4, 4'h3, 4'hc, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h5, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'h0, 4'h4, 4'h5, 4'h5, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hd, 4'hc, 4'h4, 4'h0, 4'h4, 4'hc, 4'h0, 4'h4, 4'hc, 4'hc, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h3, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h7, 4'h3, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h4, 4'hf, 4'hf, 4'hc, 4'h0, 4'hc, 4'h3, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'hc, 4'h3, 4'h3, 4'hf, 4'h1, 4'h4, 4'h3, 4'h3, 4'hf, 4'h1, 4'h5, 4'h1, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h4, 4'h1, 4'h1, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'hc, 4'hf, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'hf, 4'h5, 4'h5, 4'h0, 4'hf, 4'hd, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h1, 4'h3, 4'h1, 4'h3, 4'hc, 4'hc, 4'h5, 4'h4, 4'hf, 4'hf, 4'h0, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h5, 4'h5, 4'h3, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'hc, 4'h0, 4'h5, 4'h1, 4'h5, 4'h4, 4'h0, 4'hc, 4'hc, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h5, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'hc, 4'hc, 4'h1, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h7, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'h3, 4'hd, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h5, 4'h3, 4'hc };
assign dw_0[42] = dw_0_42[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_43 = { 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h4, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'h1, 4'h4, 4'h1, 4'h5, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'h4, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h5, 4'hc, 4'h1, 4'h4, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h1, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'hc, 4'h3, 4'hc, 4'h3, 4'hc, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'h3, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h1, 4'h1, 4'h5, 4'h1, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h4, 4'h5, 4'h4, 4'h4, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h3, 4'hc, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'hf, 4'hf, 4'h3, 4'h1, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h4, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'hc, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0 };
assign dw_0[43] = dw_0_43[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_44 = { 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h4, 4'h0, 4'hf, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h3, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hd, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h1, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hd, 4'h0, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'hc, 4'h1, 4'hc, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h7, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'hf, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'h4, 4'h4, 4'h1, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'hc, 4'hc, 4'h3, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h1, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hd, 4'h4, 4'h5, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h4, 4'h4, 4'h3, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h1, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc };
assign dw_0[44] = dw_0_44[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_45 = { 4'h5, 4'h3, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'h3, 4'h3, 4'h0, 4'hf, 4'h3, 4'hf, 4'hc, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h1, 4'h1, 4'h4, 4'h4, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h4, 4'h1, 4'h5, 4'h0, 4'h4, 4'h0, 4'h1, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'hc, 4'h3, 4'h0, 4'hf, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h1, 4'h4, 4'hc, 4'h0, 4'h3, 4'hf, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h5, 4'h4, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h5, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h1, 4'h5, 4'h1, 4'h1, 4'h5, 4'h4, 4'h4, 4'hf, 4'hc, 4'h3, 4'hc, 4'hc, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h5, 4'h1, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf };
assign dw_0[45] = dw_0_45[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_46 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[46] = dw_0_46[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_47 = { 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h3, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h5, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'h0, 4'hc, 4'h3, 4'hc, 4'hf, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'hc, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hc, 4'h3, 4'hc, 4'h5, 4'h4, 4'h5, 4'h0, 4'h5, 4'h4, 4'h5, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hc, 4'h1, 4'h4, 4'hc, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h5, 4'h4, 4'h1, 4'h4, 4'h5, 4'h1, 4'h4, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'h4, 4'h1, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'hc, 4'h3, 4'h3, 4'hf, 4'hf, 4'hc, 4'h5, 4'h7, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'hc, 4'hf, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h4, 4'hc, 4'h0, 4'h4, 4'h1, 4'h0, 4'h5, 4'h1, 4'hc, 4'hc, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h1, 4'h1, 4'h5, 4'h4, 4'h0, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'h3, 4'h3, 4'h3, 4'h3, 4'h3, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'h1, 4'h3, 4'h4, 4'h3, 4'hc, 4'h0, 4'hf, 4'h3, 4'h3, 4'h3, 4'hc, 4'h1, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h3, 4'h3, 4'hf, 4'h3, 4'hc, 4'hf, 4'h3, 4'hf, 4'h3, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf };
assign dw_0[47] = dw_0_47[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_48 = { 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h5, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h3, 4'h0, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'h5, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h1, 4'h7, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h4, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hc, 4'hf, 4'h1, 4'h3, 4'h4, 4'h4, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h5, 4'h0, 4'h1, 4'h4, 4'h5, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h1, 4'h5, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'h3, 4'h3, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h5, 4'h4, 4'h5, 4'h1, 4'h1, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h1, 4'h1, 4'h7, 4'h1, 4'h4, 4'h1, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'h1, 4'hf, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hc, 4'h3, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1 };
assign dw_0[48] = dw_0_48[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_49 = { 4'h5, 4'h4, 4'h3, 4'hf, 4'hf, 4'h0, 4'h1, 4'h5, 4'h1, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h3, 4'hf, 4'hf, 4'hf, 4'hd, 4'h5, 4'h5, 4'h5, 4'h0, 4'h7, 4'hc, 4'h4, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h5, 4'h3, 4'h5, 4'hf, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hf, 4'h5, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h5, 4'h5, 4'h0, 4'h3, 4'hf, 4'h0, 4'h1, 4'h5, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h5, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hd, 4'h5, 4'h1, 4'h5, 4'h5, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h1, 4'h4, 4'h4, 4'h4, 4'h0, 4'hc, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hd, 4'h1, 4'h5, 4'h1, 4'h5, 4'h4, 4'h0, 4'h3, 4'hc, 4'hc, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'hd, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'hf, 4'hc, 4'h3, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'hd, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h4, 4'h7, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'h5, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h4, 4'h5, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h5, 4'hf, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'hf, 4'hd, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h7, 4'h5, 4'h0, 4'h5, 4'h0, 4'h1, 4'h3, 4'h0, 4'h7, 4'h3, 4'hf, 4'hf, 4'h3, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h4, 4'h5, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h5, 4'h4, 4'h1, 4'h1, 4'h0, 4'h4, 4'h1, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hd, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h3 };
assign dw_0[49] = dw_0_49[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_50 = { 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'hc, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3, 4'hd, 4'h3, 4'h0, 4'h1, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h3, 4'hc, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'hd, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hc, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'h1, 4'h4, 4'h0, 4'hc, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h3, 4'hc, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h5, 4'h4, 4'h1, 4'h1, 4'h5, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h5, 4'h1, 4'h4, 4'h1, 4'h1, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h3, 4'hc, 4'h3, 4'hc, 4'hf, 4'h3, 4'h0, 4'hc, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'hc, 4'hf, 4'hf, 4'hc, 4'h3, 4'h1, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h4, 4'h1, 4'h1, 4'hc, 4'hf, 4'hc, 4'h3, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h1, 4'h0, 4'h1, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'hf, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h5, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'hf, 4'hc, 4'hc, 4'h0, 4'h3 };
assign dw_0[50] = dw_0_50[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_51 = { 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h3, 4'h5, 4'h4, 4'h4, 4'h4, 4'h5, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h1, 4'h4, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h1, 4'h5, 4'h5, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'h5, 4'hc, 4'hc, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'h3, 4'hf, 4'h5, 4'h5, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'hf, 4'hf, 4'h1, 4'h3, 4'h3, 4'h0, 4'hf, 4'hd, 4'h5, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'h0, 4'h5, 4'hc, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'h1, 4'hc, 4'h1, 4'h5, 4'h5, 4'h1, 4'h0, 4'h5, 4'h7, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'hc, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h4, 4'h1, 4'h4, 4'h1, 4'h4, 4'h5, 4'h1, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h7, 4'h0, 4'h3, 4'hd, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h4, 4'h4, 4'h0, 4'hc, 4'hd, 4'h5, 4'h4, 4'hf, 4'hf, 4'h0, 4'hc, 4'hf, 4'h0, 4'h3, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h3, 4'hf, 4'hc, 4'h3, 4'h4, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'h0, 4'h3, 4'hf, 4'h0, 4'hf, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h4, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'h4, 4'h5, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'hf, 4'h3, 4'h3, 4'h3, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h0, 4'h0, 4'h4, 4'hf, 4'h3, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hd, 4'h4, 4'h5, 4'h0, 4'hf, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h4, 4'hc, 4'hc, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'hc, 4'hf, 4'h0, 4'h3, 4'hf, 4'hc, 4'hc, 4'hc, 4'hc, 4'hf, 4'hf, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hd, 4'h0, 4'h3, 4'hc, 4'hf, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd };
assign dw_0[51] = dw_0_51[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_52 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'h3, 4'hc, 4'h3, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hf, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h5, 4'h4, 4'h1, 4'h1, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h0, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'h5, 4'h1, 4'h0, 4'h3, 4'hf, 4'h0, 4'h3, 4'h3, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'hc, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'h5, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h1, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h4, 4'h1, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'hc, 4'h0, 4'h1, 4'h3, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'hc, 4'h3, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[52] = dw_0_52[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_53 = { 4'hf, 4'hf, 4'h0, 4'h5, 4'h0, 4'h5, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h1, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'hf, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h1, 4'h0, 4'h4, 4'h5, 4'h1, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'hf, 4'h3, 4'hc, 4'hc, 4'hc, 4'hc, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'hf, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h4, 4'h3, 4'h0, 4'hc, 4'h1, 4'h1, 4'hc, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h4, 4'h5, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'h3, 4'hf, 4'h1, 4'h4, 4'hc, 4'hd, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'h3, 4'hf, 4'hc, 4'hd, 4'hd, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'h3, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h3, 4'hf, 4'h5, 4'h1, 4'h1, 4'h1, 4'h1, 4'h1, 4'h4, 4'h4, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h4, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h5, 4'h0, 4'h7, 4'hf, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h5, 4'h7, 4'h5, 4'h1, 4'h1, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h1, 4'h0, 4'h7, 4'h5, 4'h0, 4'h5, 4'h5, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hc, 4'hc, 4'h3, 4'h3, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'h0, 4'h3, 4'h4, 4'h1, 4'h3, 4'h0, 4'hd, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5 };
assign dw_0[53] = dw_0_53[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_54 = { 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h0, 4'h5, 4'h4, 4'h4, 4'h5, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h1, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h3, 4'hc, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hf, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'hd, 4'h1, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h1, 4'h0, 4'h4, 4'h4, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h1, 4'h5, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'hf };
assign dw_0[54] = dw_0_54[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_55 = { 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hc, 4'hf, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'h4, 4'hc, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'h4, 4'h5, 4'h4, 4'h5, 4'h0, 4'h5, 4'h4, 4'h5, 4'h3, 4'h3, 4'h3, 4'hf, 4'hf, 4'h3, 4'h0, 4'hd, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'h0, 4'h3, 4'h4, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h4, 4'h5, 4'h4, 4'h0, 4'h5, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h1, 4'h4, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h4, 4'h3, 4'hc, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h4, 4'h4, 4'h5, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'h0, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'hc, 4'hf, 4'hc, 4'h3, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h0, 4'h4, 4'h4, 4'h5, 4'h4, 4'h0, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h5, 4'h4, 4'h4, 4'h1, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'h1, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h7, 4'hc, 4'hf, 4'h3, 4'h0, 4'h3, 4'h3, 4'h3, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h7, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hc, 4'h3, 4'hc, 4'h3, 4'hf, 4'hc, 4'hc, 4'hf, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1 };
assign dw_0[55] = dw_0_55[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_56 = { 4'h3, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h3, 4'h0, 4'h3, 4'hc, 4'h1, 4'h4, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h0, 4'h4, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'h7, 4'hf, 4'h3, 4'h4, 4'h1, 4'h1, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'h4, 4'h5, 4'h1, 4'h5, 4'h7, 4'h0, 4'h5, 4'h5, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'hf, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h5, 4'h0, 4'hc, 4'h4, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h1, 4'h5, 4'h1, 4'h0, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h1, 4'hc, 4'h0, 4'h4, 4'h0, 4'hf, 4'hc, 4'h3, 4'hf, 4'h4, 4'h1, 4'h5, 4'h0, 4'h4, 4'h4, 4'h5, 4'h5, 4'h3, 4'h3, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h3, 4'h3, 4'h3, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h3, 4'h1, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h3, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'hf, 4'h0, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h4, 4'h1, 4'h4, 4'h5, 4'h0, 4'h1, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'hf, 4'h3, 4'h3, 4'hc, 4'hf, 4'hf, 4'hd, 4'hf, 4'hf, 4'h0, 4'hc, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4, 4'h0, 4'hd, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'h1, 4'h5, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0 };
assign dw_0[56] = dw_0_56[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_57 = { 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'h3, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'hf, 4'h0, 4'hf, 4'h0, 4'h5, 4'h1, 4'h1, 4'h5, 4'h1, 4'h5, 4'h1, 4'h4, 4'h7, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'h5, 4'h0, 4'h1, 4'h1, 4'h1, 4'h0, 4'h1, 4'hf, 4'hf, 4'h0, 4'h7, 4'h3, 4'h5, 4'hf, 4'h3, 4'h5, 4'h5, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'hc, 4'h0, 4'hf, 4'h3, 4'hc, 4'hf, 4'h0, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'h0, 4'hf, 4'hf, 4'hc, 4'hf, 4'h1, 4'h5, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h7, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'h1, 4'h4, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'hc, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'hc, 4'h4, 4'h3, 4'hf, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'hc, 4'h3, 4'hf, 4'hc, 4'h0, 4'h3, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'hc, 4'hc, 4'h1, 4'hc, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'hf, 4'h1, 4'h0, 4'h4, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h7, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h3, 4'h5, 4'hc, 4'hc, 4'h0, 4'hc, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hd, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'hf, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'hc, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h5, 4'h4, 4'h1, 4'h1, 4'h5, 4'h0, 4'h5, 4'h5, 4'hd, 4'hf, 4'h3, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h3, 4'hc, 4'hf, 4'h1, 4'h0, 4'hf, 4'hc, 4'hf, 4'h3, 4'hc, 4'hf, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hd, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h7, 4'hc, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'hd };
assign dw_0[57] = dw_0_57[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_58 = { 4'hf, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'hc, 4'hc, 4'hc, 4'h0, 4'hf, 4'hf, 4'h7, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hd, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h3, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'hf, 4'h3, 4'h3, 4'hc, 4'h0, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'hc, 4'h3, 4'hf, 4'hc, 4'h1, 4'h5, 4'hf, 4'hc, 4'h1, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h5, 4'h1, 4'h0, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'hd, 4'h5, 4'h5, 4'h3, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h5, 4'h4, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h1, 4'h5, 4'h4, 4'h0, 4'hf, 4'hf, 4'h0, 4'h1, 4'h5, 4'h7, 4'h0, 4'hf, 4'hc, 4'hf, 4'h3, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'hf, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h3, 4'hc, 4'h3, 4'hc, 4'hf, 4'h3, 4'h1, 4'h0, 4'h4, 4'h4, 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h5, 4'h3, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h4, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h1, 4'h5, 4'h5, 4'h1, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'hc, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hd, 4'h3, 4'h0, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'hf, 4'hf, 4'hc, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'h3, 4'h0, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h1 };
assign dw_0[58] = dw_0_58[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_59 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[59] = dw_0_59[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_60 = { 4'h3, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'h1, 4'h3, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'h4, 4'h1, 4'h1, 4'h5, 4'h1, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'hc, 4'hc, 4'h4, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h1, 4'h1, 4'h5, 4'h4, 4'hd, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h0, 4'h5, 4'h5, 4'hf, 4'hc, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h5, 4'h4, 4'h4, 4'h4, 4'h1, 4'h1, 4'h5, 4'h4, 4'h1, 4'h1, 4'h4, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h4, 4'h3, 4'h3, 4'hc, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'h1, 4'hf, 4'hc, 4'h0, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'h3, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h5, 4'h1, 4'h5, 4'hc, 4'hc, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h4, 4'h0, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h5, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h4, 4'h4, 4'h5, 4'h4, 4'h4, 4'h5, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hc, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'h1, 4'h3, 4'hc, 4'hd, 4'h3, 4'hf, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h4, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h3, 4'h1, 4'hf, 4'h1, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'hf, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h5, 4'h4, 4'h4, 4'h1, 4'h0, 4'h4, 4'h5, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h4, 4'h4, 4'h0 };
assign dw_0[60] = dw_0_60[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_61 = { 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'hc, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h5, 4'h1, 4'h7, 4'h5, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'hf, 4'hf, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h1, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'hd, 4'h3, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h1, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'hf, 4'h3, 4'h3, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h4, 4'h4, 4'h1, 4'h1, 4'h4, 4'h0, 4'h5, 4'h0, 4'h1, 4'h4, 4'h1, 4'h7, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'hc, 4'h4, 4'h4, 4'hc, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h3, 4'hc, 4'hc, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h4, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h3, 4'hf, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h1, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h7, 4'h5, 4'h1, 4'h4, 4'h5, 4'h0, 4'h1, 4'h5, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'hc, 4'hd, 4'h5, 4'h1, 4'h5, 4'h0, 4'h5, 4'h4, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hd, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5 };
assign dw_0[61] = dw_0_61[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_62 = { 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h1, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'hf, 4'h0, 4'hf, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h3, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'h5, 4'h0, 4'h5, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h1, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h0, 4'h5, 4'h4, 4'h4, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'h0, 4'hc, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h7, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hd, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hd, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h5, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h1, 4'h4 };
assign dw_0[62] = dw_0_62[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_63 = { 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h1, 4'h4, 4'h3, 4'hc, 4'h3, 4'hf, 4'h0, 4'h3, 4'hc, 4'h3, 4'h1, 4'h4, 4'h0, 4'h3, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h3, 4'h5, 4'h5, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h5, 4'h0, 4'h4, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h3, 4'hc, 4'h0, 4'hc, 4'h7, 4'h0, 4'h3, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h3, 4'h0, 4'h0, 4'hf, 4'hc, 4'h7, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'h5, 4'hc, 4'h1, 4'h4, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'hd, 4'h5, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h5, 4'h4, 4'h5, 4'h1, 4'h1, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h1, 4'h1, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'h0, 4'hc, 4'hf, 4'hc, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h4, 4'h5, 4'h4, 4'h1, 4'h1, 4'h1, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'h3, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'hf, 4'h4, 4'hc, 4'h1, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h4, 4'h5, 4'h4, 4'h0, 4'h4, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h1, 4'h4, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'h0, 4'h5, 4'h4, 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h4, 4'h1, 4'h4, 4'h5, 4'h4, 4'h1, 4'h0, 4'h4, 4'h5, 4'h4, 4'h4, 4'hc, 4'h4, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3 };
assign dw_0[63] = dw_0_63[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_64 = { 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'hf, 4'h1, 4'h4, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h5, 4'hd, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'h3, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'h3, 4'h3, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'h0, 4'h3, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h3, 4'hf, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h3, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hf, 4'h1, 4'h3, 4'hf, 4'h3, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h4, 4'h5, 4'h1, 4'h4, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'hf, 4'h3, 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[64] = dw_0_64[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_65 = { 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h3, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h4, 4'h1, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h3, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h5, 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'h3, 4'h0, 4'h4, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h1, 4'h5, 4'h4, 4'h1, 4'h4, 4'h0, 4'hc, 4'hc, 4'h3, 4'hf, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'hf, 4'h3, 4'h3, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'hf, 4'hc, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'hf, 4'h3, 4'h3, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0 };
assign dw_0[65] = dw_0_65[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_66 = { 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h3, 4'hf, 4'h0, 4'hc, 4'h1, 4'h3, 4'h3, 4'h0, 4'h4, 4'h1, 4'h5, 4'h0, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h5, 4'hc, 4'hc, 4'hc, 4'hc, 4'hf, 4'h0, 4'hc, 4'h3, 4'h3, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'h1, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'h0, 4'h1, 4'h3, 4'hc, 4'hd, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'hf, 4'h3, 4'h0, 4'h3, 4'hc, 4'hf, 4'h3, 4'hf, 4'hc, 4'hc, 4'hd, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hd, 4'h5, 4'h4, 4'h1, 4'h4, 4'h1, 4'h4, 4'h0, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hc, 4'hd, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'hf, 4'hc, 4'hc, 4'hc, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'hf, 4'h4, 4'h4, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h4, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h7, 4'hc, 4'h3, 4'h3, 4'h3, 4'h0, 4'hf, 4'hf, 4'h3, 4'h3, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h4, 4'h4, 4'h4, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h5, 4'h1, 4'h4, 4'h0, 4'h7, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h7, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'h4, 4'h3, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h4, 4'h4, 4'h1, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'hf, 4'h1, 4'hc, 4'h7, 4'hc, 4'hc, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5 };
assign dw_0[66] = dw_0_66[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_67 = { 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h4, 4'hd, 4'h1, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h0, 4'h1, 4'h5, 4'h1, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'hf, 4'hc, 4'hf, 4'hc, 4'hf, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h3, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h4, 4'h1, 4'h1, 4'h5, 4'h1, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h1, 4'h4, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h4, 4'h5, 4'h0, 4'h1, 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h5, 4'h4, 4'h5, 4'h1, 4'h4, 4'h5, 4'h4, 4'hf, 4'hf, 4'h0, 4'hc, 4'hc, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h5, 4'h0, 4'h4, 4'h1, 4'h5, 4'h1, 4'h5, 4'h4, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'hc, 4'hf, 4'hc, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'hc, 4'h5, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h3, 4'h0, 4'h4, 4'h5, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'h0, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'h0, 4'h5, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h1, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h1, 4'h7, 4'h3, 4'h4, 4'hf, 4'h1, 4'h7, 4'h0 };
assign dw_0[67] = dw_0_67[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_68 = { 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'hf, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h4, 4'h4, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'hf, 4'h3, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h7, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h4, 4'h5, 4'h1, 4'h1, 4'h1, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'hf, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'h5, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'hc, 4'h3, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'hc, 4'hf, 4'h3, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'hd, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'h3, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h5, 4'h4, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'hc, 4'hc, 4'hc, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0 };
assign dw_0[68] = dw_0_68[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_69 = { 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h1, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h4, 4'h1, 4'h5, 4'h4, 4'h5, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'hd, 4'h5, 4'h0, 4'h1, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h4, 4'h4, 4'hc, 4'h4, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h3, 4'h4, 4'hc, 4'h0, 4'h5, 4'h1, 4'h4, 4'h1, 4'h4, 4'hc, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h5, 4'hf, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hd, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hc, 4'hf, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'h3, 4'h3, 4'hc, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h1, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'h3, 4'h3, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'hd, 4'h7, 4'hc, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h0, 4'hc, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h1, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h5, 4'h5, 4'h4, 4'h1, 4'h4, 4'h1, 4'h0, 4'h1, 4'h5, 4'h5, 4'h1, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h1, 4'h0, 4'h1, 4'hf, 4'h3, 4'h0, 4'h3, 4'h3, 4'hc, 4'h1, 4'h1, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'h5, 4'h3, 4'h4, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h5, 4'h1 };
assign dw_0[69] = dw_0_69[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_70 = { 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hd, 4'hc, 4'h0, 4'h4, 4'h7, 4'h3, 4'hc, 4'h3, 4'h3, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'hd, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h0, 4'h5, 4'h4, 4'h1, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h1, 4'h0, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'hc, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4, 4'h4, 4'hc, 4'h4, 4'h4, 4'h0, 4'h1, 4'hc, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'h3, 4'hf, 4'h4, 4'h0, 4'h1, 4'h0, 4'h5, 4'h5, 4'h1, 4'h0, 4'h4, 4'h1, 4'h5, 4'h1, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h3, 4'hd, 4'h3, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'hf, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h4, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h7, 4'h3, 4'hf, 4'h0, 4'hf, 4'hc, 4'h1, 4'h4, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5, 4'h1, 4'h4, 4'h5, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'h3, 4'h3, 4'h0 };
assign dw_0[70] = dw_0_70[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_71 = { 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h1, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'hc, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h1, 4'h5, 4'h4, 4'h1, 4'h0, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'hf, 4'h3, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hf, 4'hc, 4'h3, 4'hf, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h0, 4'h4, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h5, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h0, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h0, 4'h5, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h4, 4'h1, 4'h5, 4'h5, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0 };
assign dw_0[71] = dw_0_71[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_72 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[72] = dw_0_72[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_73 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'hf, 4'h3, 4'hc, 4'h3, 4'hd, 4'h3, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h1, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[73] = dw_0_73[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_74 = { 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1 };
assign dw_0[74] = dw_0_74[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_75 = { 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'hc, 4'hc, 4'hf, 4'h3, 4'h3, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h1, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h3, 4'hc, 4'h3, 4'hf, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h5, 4'h4, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'h0, 4'h1, 4'h5, 4'h1, 4'h0, 4'h1, 4'h5, 4'h1, 4'h5, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'hc, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'h4, 4'h5, 4'h3, 4'h3, 4'hf, 4'h0, 4'hf, 4'hf, 4'h3, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'h1, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'h1, 4'h0 };
assign dw_0[75] = dw_0_75[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_76 = { 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h3, 4'hf, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'hc, 4'hf, 4'hf, 4'h3, 4'h3, 4'hf, 4'hc, 4'hf, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h4, 4'hf, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'hc, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'hf, 4'hf, 4'h0, 4'h3, 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h5, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h0, 4'h5, 4'h1, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'hf, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3 };
assign dw_0[76] = dw_0_76[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_77 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h4, 4'h4, 4'h5, 4'h1, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'hc, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h5, 4'h1, 4'h4, 4'h4, 4'h1, 4'h1, 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'h3, 4'h3, 4'hc, 4'hf };
assign dw_0[77] = dw_0_77[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_78 = { 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h7, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'h0, 4'h1, 4'h1, 4'h0, 4'h4, 4'hd, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h1, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'h3, 4'h3, 4'hc, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h1, 4'h3, 4'h0, 4'hd, 4'h0, 4'h0, 4'hc, 4'h1, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'h5, 4'h4, 4'h5, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf };
assign dw_0[78] = dw_0_78[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_79 = { 4'h5, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h5, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'h4, 4'h5, 4'h4, 4'h5, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'hf, 4'hc, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'hf, 4'h4, 4'h5, 4'h5, 4'h4, 4'h1, 4'h1, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h1, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'h1, 4'h5, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'hf, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h4, 4'h4, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'h3, 4'h3, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h5, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hc, 4'h3, 4'hf, 4'hf, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0 };
assign dw_0[79] = dw_0_79[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_80 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[80] = dw_0_80[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_81 = { 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h0, 4'h1, 4'h1, 4'h0, 4'h4, 4'h1, 4'h4, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'hf, 4'h3, 4'h3, 4'hf, 4'h4, 4'h0, 4'h4, 4'h5, 4'h4, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'hc, 4'h3, 4'h1, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h3, 4'hf, 4'h0, 4'hc, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'h0, 4'h4, 4'hd, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'h5, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'hd, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h1, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'h4, 4'hd, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'h4, 4'h7, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'h1, 4'h5, 4'h4, 4'h1, 4'h5, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h4, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h4, 4'h4, 4'hc, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h7, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'h0, 4'h1, 4'h1, 4'h5, 4'h0, 4'hc, 4'h4, 4'h1, 4'h5, 4'h4, 4'h1, 4'h3, 4'h1, 4'h0, 4'h3, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h0, 4'h1, 4'h5, 4'h0, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h1, 4'h4, 4'h7, 4'h1, 4'h0, 4'h1, 4'h0, 4'hf, 4'h4, 4'h0, 4'h5, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'h1, 4'h0, 4'h5, 4'h0, 4'h1, 4'h1, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'h4, 4'h0, 4'hc, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h4, 4'h1, 4'h1, 4'h1, 4'h5, 4'h3, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0 };
assign dw_0[81] = dw_0_81[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_82 = { 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'hc, 4'hc, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'h3, 4'h3, 4'h3, 4'h0, 4'hf, 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'h4, 4'h1, 4'h0, 4'h5, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'hc, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h3, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h4, 4'h1, 4'h1, 4'h4, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h4, 4'h5, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'h3, 4'h3, 4'hf, 4'hc, 4'hf, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h1, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'hc, 4'h5, 4'h0, 4'h3, 4'h1, 4'hc, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'hc, 4'h3, 4'h3, 4'h3, 4'hc, 4'h3, 4'hc, 4'hc, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'hf, 4'hf, 4'h3, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h1, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h7, 4'h0, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hd, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hd, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'hf, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'h0, 4'hc };
assign dw_0[82] = dw_0_82[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_83 = { 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hd, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'hc, 4'hf, 4'h3, 4'h3, 4'h3, 4'hf, 4'hf, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'hc, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'h3, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hd, 4'h4, 4'h4, 4'h4, 4'h0, 4'h1, 4'h1, 4'h3, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'hc, 4'h3, 4'h5, 4'h5, 4'h1, 4'h0, 4'h5, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'hc, 4'hf, 4'hc, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h3, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h4, 4'h4, 4'h1, 4'h4, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h5, 4'h1, 4'h1, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h5, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h4, 4'h1, 4'h1, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h4, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h1, 4'h5, 4'hf, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h1, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'hf, 4'hc, 4'hc, 4'hd, 4'h0, 4'h4, 4'h0, 4'h5, 4'h1, 4'h1, 4'h7 };
assign dw_0[83] = dw_0_83[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_84 = { 4'h3, 4'hc, 4'hc, 4'hc, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'h3, 4'hf, 4'h3, 4'hc, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h5, 4'h1, 4'h0, 4'h4, 4'h3, 4'h3, 4'hf, 4'hc, 4'hf, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h5, 4'h5, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[84] = dw_0_84[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_85 = { 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h5, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hc, 4'h3, 4'hf, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h3, 4'h3, 4'h3, 4'h3, 4'hd, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h3, 4'h3, 4'hc, 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'h5, 4'h4, 4'h1, 4'h1, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h1, 4'h5, 4'h4, 4'h1, 4'h1, 4'h1, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h5, 4'h0, 4'h5, 4'h1, 4'h4, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h4, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h5, 4'h1, 4'h1, 4'h1, 4'h4, 4'h5, 4'h4, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h5, 4'h0, 4'hf, 4'hf, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'h1, 4'h4, 4'h5, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h1, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h5, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h1, 4'h1, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h4, 4'hf, 4'h3, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc };
assign dw_0[85] = dw_0_85[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_86 = { 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h4, 4'h1, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'hc, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h5, 4'h4, 4'h0, 4'h1, 4'h5, 4'h4, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h1, 4'h5, 4'h1, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h3, 4'h3, 4'hf, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h5, 4'h4, 4'hc, 4'h0, 4'h5, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'hf, 4'h3, 4'hc, 4'h3, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h1, 4'h1, 4'h4, 4'hd, 4'h4, 4'h4, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'hf, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h1, 4'h3, 4'h0, 4'h4, 4'hd, 4'h5, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'h5, 4'h5, 4'h1, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h1, 4'h1, 4'h0, 4'h1, 4'h5, 4'h5, 4'h0, 4'h4, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1 };
assign dw_0[86] = dw_0_86[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_87 = { 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'h1, 4'h5, 4'h1, 4'h5, 4'h4, 4'h0, 4'h5, 4'h1, 4'hf, 4'hc, 4'h1, 4'h1, 4'h0, 4'h3, 4'hc, 4'hf, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h4, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h4, 4'hc, 4'hc, 4'hc, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h1, 4'h5, 4'h4, 4'h0, 4'hc, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hf, 4'h3, 4'h5, 4'h5, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'hc, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'hf, 4'hc, 4'hc, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h4, 4'h1, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc };
assign dw_0[87] = dw_0_87[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_88 = { 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h1, 4'h1, 4'h5, 4'hd, 4'h0, 4'h0, 4'h7, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h1, 4'hd, 4'h4, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h4, 4'h1, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hc, 4'h0, 4'h5, 4'h0, 4'h4, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hd, 4'h4, 4'h1, 4'h5, 4'h5, 4'h4, 4'hd, 4'h0, 4'h1, 4'h4, 4'h1, 4'h5, 4'h0, 4'h1, 4'h5, 4'h1, 4'h0, 4'h1, 4'h3, 4'hf, 4'hc, 4'h3, 4'h3, 4'h3, 4'hf, 4'h7, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h1, 4'h1, 4'h0, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h7, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'hf, 4'h0, 4'hf, 4'h3, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3, 4'h5, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'h5, 4'h1, 4'h4, 4'h5, 4'h1, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'h0, 4'hc, 4'h3, 4'hf, 4'hc, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'h4, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'hd, 4'h0, 4'h5, 4'h1, 4'h5, 4'h0, 4'h5, 4'h1, 4'h4, 4'h0, 4'hf, 4'h1, 4'h0, 4'h1, 4'h3, 4'hf, 4'h3, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'hd, 4'h4, 4'h1, 4'h0, 4'h5, 4'h5, 4'hd, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h5, 4'h1, 4'h1, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'hf, 4'hc, 4'hc, 4'h3, 4'hf, 4'h3, 4'hc, 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'hf, 4'hf, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h3, 4'hc, 4'hf, 4'h3, 4'hf, 4'h3, 4'hf, 4'hd, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'hf, 4'h0, 4'h3, 4'hf, 4'h0, 4'hd, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h5, 4'h0, 4'h5, 4'hf, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'h1, 4'hc, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h7, 4'hd, 4'hc, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5 };
assign dw_0[88] = dw_0_88[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_89 = { 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h5, 4'h1, 4'h1, 4'h4, 4'h0, 4'hf, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h5, 4'h1, 4'h4, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h5, 4'h4, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h1, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3 };
assign dw_0[89] = dw_0_89[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_90 = { 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h4, 4'h5, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h7, 4'h1, 4'h4, 4'h1, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hd, 4'h4, 4'hc, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'h5, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h7, 4'h0, 4'h4, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h5, 4'h4, 4'h0, 4'h4, 4'h5, 4'h0, 4'h3, 4'h3, 4'hc, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h7, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'hc, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'h3, 4'h4, 4'hc, 4'h0, 4'hf, 4'h4, 4'h4, 4'h4, 4'h1, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h5, 4'h0, 4'h4, 4'h4, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h4, 4'h0, 4'h4, 4'h5, 4'h1, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h5, 4'h4, 4'h5, 4'h1, 4'hc, 4'h1, 4'h3, 4'h3, 4'hf, 4'hc, 4'h7, 4'h0, 4'h0, 4'hd, 4'h5, 4'h5, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'hc, 4'h0, 4'h4, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'hd, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3, 4'h4, 4'hf, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h3, 4'h3, 4'h5, 4'hc, 4'h4, 4'h4, 4'h5, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h0, 4'h1, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'h7, 4'h1, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h7, 4'h1, 4'h5, 4'h1, 4'h4, 4'h4, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h5, 4'h3, 4'h3, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'hf, 4'hc, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h7, 4'h0, 4'hc, 4'h3, 4'hf, 4'h0, 4'h1, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h5, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0 };
assign dw_0[90] = dw_0_90[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_91 = { 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'h0, 4'h3, 4'hd, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h4, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h7, 4'h4, 4'h1, 4'h3, 4'h5, 4'h1, 4'h0, 4'hd, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'hc, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'h3, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'hc, 4'hf, 4'hc, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h1, 4'h4, 4'h0, 4'h1, 4'h1, 4'h5, 4'hc, 4'h5, 4'h5, 4'h1, 4'hf, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h1, 4'hf, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h4, 4'h3, 4'hc, 4'hc, 4'hc, 4'hf, 4'h3, 4'h5, 4'h4, 4'h1, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h0, 4'h5, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'hc, 4'h3, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h5, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h3, 4'hf, 4'h1, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h5, 4'h5, 4'h7, 4'h5, 4'h5, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'hf, 4'h0, 4'h3, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h7, 4'hc, 4'hc, 4'h0, 4'hc, 4'h1, 4'h3, 4'h7, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h1, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h1, 4'h0, 4'hf, 4'hc, 4'hf, 4'h7, 4'h4, 4'h5, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h3, 4'h4, 4'h1, 4'h4, 4'h1, 4'h1, 4'h5, 4'h5, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h7, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'hd, 4'h3, 4'h3, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h1 };
assign dw_0[91] = dw_0_91[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_92 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h0, 4'h5, 4'h4, 4'h0, 4'h3, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'hf, 4'h0, 4'hc, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h1, 4'hf, 4'hc, 4'h4, 4'h1, 4'h5, 4'h0, 4'h3, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'hf, 4'hf, 4'h0, 4'h7, 4'h0, 4'h5, 4'hf, 4'h3, 4'h5, 4'h3, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h4, 4'h4, 4'hf, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h1, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h1, 4'h0, 4'h1, 4'h5, 4'h0, 4'hd, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h4, 4'h1, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hf, 4'h5, 4'h4, 4'h1, 4'h4, 4'hd, 4'h7, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'h0, 4'h5, 4'h0, 4'hc, 4'h4, 4'h0, 4'hf, 4'hc, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h1, 4'h4, 4'hf, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'hc, 4'h3, 4'h0, 4'h1, 4'h5, 4'h3, 4'hf, 4'h3, 4'h1, 4'h3, 4'h0, 4'h3, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h4, 4'h0, 4'h1, 4'h0, 4'h5, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'hc, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'h5, 4'h3, 4'h1, 4'h1, 4'h1, 4'h5, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'h5, 4'h3, 4'hc, 4'h5, 4'hf, 4'h4, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'h0, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h1, 4'h1, 4'h1, 4'h4, 4'h4, 4'h0, 4'hc, 4'h4, 4'h1, 4'h4, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'h0, 4'h5, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'hf, 4'h1, 4'hf, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h1, 4'h3, 4'h3, 4'h3, 4'hc, 4'h1, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h1, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h4, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h7, 4'h0, 4'hd, 4'h4, 4'hc, 4'h0, 4'h0, 4'h1, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'hd, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'h1, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'hf, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'hc, 4'h0, 4'h7, 4'h7, 4'hc, 4'h0, 4'hf, 4'hf, 4'hc, 4'h3, 4'hd };
assign dw_0[92] = dw_0_92[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_93 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[93] = dw_0_93[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_94 = { 4'h4, 4'h1, 4'h4, 4'h4, 4'h1, 4'h4, 4'h4, 4'h0, 4'hf, 4'hc, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0, 4'h3, 4'hf, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h5, 4'h7, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'hc, 4'h4, 4'h7, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'hc, 4'h0, 4'h5, 4'h4, 4'h4, 4'h5, 4'h0, 4'hf, 4'h1, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'hd, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h7, 4'h4, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'h1, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'hd, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'hf, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h0, 4'h5, 4'h0, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'hc, 4'h0, 4'h5, 4'hf, 4'h0, 4'h4, 4'h3, 4'h3, 4'hc, 4'h0, 4'h3, 4'h4, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'h3, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h5, 4'h5, 4'h3, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hd, 4'hc, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'hd, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h1, 4'h5, 4'h4, 4'hf, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'hc, 4'h3, 4'hc, 4'h4, 4'h0, 4'h1, 4'hf, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h4, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd };
assign dw_0[94] = dw_0_94[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_95 = { 4'h0, 4'h3, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'hf, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[95] = dw_0_95[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_96 = { 4'h1, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h1, 4'h5, 4'h4, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h4, 4'h4, 4'h0, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3 };
assign dw_0[96] = dw_0_96[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_97 = { 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'h5, 4'h1, 4'h4, 4'h4, 4'h1, 4'h4, 4'h5, 4'h5, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hd, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h3, 4'h3, 4'h7, 4'h3, 4'hf, 4'hc, 4'hc, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'hc, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h1, 4'h1, 4'h1, 4'h5, 4'h5, 4'h7, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'h5, 4'h1, 4'h4, 4'h5, 4'h4, 4'h5, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'h3, 4'h0, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h0, 4'h4, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h5, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'hc, 4'h4, 4'h7, 4'hc, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'hc, 4'h3, 4'h3, 4'hc, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h1, 4'h3, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h7, 4'h5, 4'h1, 4'h7, 4'h0, 4'h0, 4'h7, 4'hc, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'hc, 4'h3, 4'h0, 4'h1, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf };
assign dw_0[97] = dw_0_97[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_98 = { 4'hf, 4'h0, 4'hc, 4'h0, 4'hf, 4'h3, 4'h3, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h5, 4'h1, 4'h5, 4'h1, 4'h5, 4'h0, 4'h1, 4'h4, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h7, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h1, 4'h4, 4'h1, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'h0, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h4, 4'h1, 4'h0, 4'h1, 4'h1, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h3, 4'h0, 4'h3, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5 };
assign dw_0[98] = dw_0_98[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_99 = { 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h0, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h1, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'hc, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h5, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'h1, 4'h3, 4'hf, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hc, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h1, 4'h5, 4'h4, 4'h4, 4'h4, 4'h1, 4'h1, 4'h5, 4'h0, 4'h5, 4'h0, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'hc, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h5, 4'h4, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h1, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'hc, 4'hf, 4'h3, 4'hc, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hd, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'hc, 4'hc, 4'hf, 4'hc, 4'h3, 4'hc, 4'h3, 4'hf, 4'hc, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h1, 4'h1, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc };
assign dw_0[99] = dw_0_99[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_100 = { 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h1, 4'h5, 4'h4, 4'h0, 4'h5, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h1, 4'h4, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'hc, 4'h5, 4'h4, 4'h1, 4'h1, 4'h0, 4'h4, 4'h3, 4'h5, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'hc, 4'h3, 4'hf, 4'hf, 4'h0, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3, 4'h3, 4'hc, 4'h1, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'hf, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'hc, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h5, 4'h0, 4'h4, 4'h4, 4'h4, 4'h1, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h3, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h7, 4'h0, 4'h5, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h5, 4'h0, 4'h7, 4'h0, 4'h4, 4'h4, 4'h3, 4'h0, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h4, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h1, 4'h5, 4'h1, 4'h0, 4'h4, 4'h5, 4'h1, 4'h3, 4'hc, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h4, 4'h5, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf };
assign dw_0[100] = dw_0_100[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_101 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'hc, 4'h3, 4'hc, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'hc, 4'h3, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h3, 4'h3, 4'h5, 4'h4, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hc, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h1, 4'h4, 4'h5, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'hc, 4'hf, 4'h3, 4'h3, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'h1, 4'h0, 4'h5, 4'h0, 4'hc, 4'hc, 4'h3, 4'hf, 4'hc, 4'h0, 4'h3, 4'hf, 4'hc, 4'hc, 4'h3, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h1, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hd, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'hc, 4'h3, 4'h3, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf };
assign dw_0[101] = dw_0_101[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_102 = { 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h4, 4'h1, 4'h1, 4'h5, 4'h0, 4'h1, 4'h5, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'hf, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'h1, 4'h7, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h1, 4'h0, 4'h5, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0 };
assign dw_0[102] = dw_0_102[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_103 = { 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h4, 4'h1, 4'h5, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hd, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h3, 4'hc, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'hc, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h5, 4'h0, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h1, 4'h1, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'h1, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h1, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h1, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h7, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h5, 4'h0, 4'h1, 4'h7, 4'h4, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h1, 4'h4, 4'h1, 4'h4, 4'h5, 4'h0, 4'hf, 4'hf, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h4, 4'h5, 4'h0, 4'h4, 4'h5, 4'h5, 4'h1, 4'h0, 4'h1, 4'h1, 4'h4, 4'hc, 4'hc, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h5, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h5, 4'hf, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5 };
assign dw_0[103] = dw_0_103[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_104 = { 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'h3, 4'h3, 4'h3, 4'h3, 4'hc, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h5, 4'h1, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h3, 4'h1, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hd, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h4, 4'h1, 4'h0, 4'h5, 4'h1, 4'h0, 4'h4, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hc, 4'hc, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h4, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h4, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'h5, 4'h1, 4'h5, 4'h1, 4'h1, 4'h1, 4'h1, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h1, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h0, 4'h5, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h1, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'h5, 4'h4, 4'h5, 4'h4, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hd, 4'h1, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'h0, 4'h4, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'h1, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h1, 4'hc, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'h3, 4'hf, 4'h3, 4'h3, 4'h3, 4'h3, 4'hc, 4'h3, 4'hf, 4'h3, 4'hc, 4'hf, 4'hc, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf };
assign dw_0[104] = dw_0_104[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_105 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h4, 4'h4, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5, 4'h1, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h1, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h3, 4'h3, 4'hc, 4'hf, 4'h3, 4'h3, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h0, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'h3, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hf, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h1, 4'hc, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf };
assign dw_0[105] = dw_0_105[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_106 = { 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h5, 4'h5, 4'h3, 4'hf, 4'h0, 4'h1, 4'h5, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'hf, 4'h3, 4'hc, 4'h3, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h5, 4'h0, 4'h1, 4'h4, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'hf, 4'h5, 4'h0, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h5, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h1, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h1, 4'h7, 4'hc, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h4, 4'h0, 4'h4, 4'hf, 4'h0, 4'hc, 4'hc, 4'hc, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h4, 4'h0, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'hd, 4'h1, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h4, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'h0, 4'h4, 4'h4, 4'h5, 4'h4, 4'h0, 4'h1, 4'h1, 4'h4, 4'h5, 4'h5, 4'h1, 4'h4, 4'h4, 4'h0, 4'h5, 4'h5, 4'hf, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h1, 4'h4, 4'h1, 4'h1, 4'h0, 4'hc, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h5, 4'h0, 4'h4, 4'h4, 4'h7, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h5, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h4, 4'h4, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h1, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'h3, 4'hc, 4'h3, 4'h3 };
assign dw_0[106] = dw_0_106[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_107 = { 4'h5, 4'h5, 4'h3, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'hf, 4'hc, 4'h0, 4'h4, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hc, 4'h5, 4'h5, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'hd, 4'h1, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'h4, 4'h0, 4'hf, 4'h3, 4'hc, 4'hc, 4'h0, 4'h5, 4'h0, 4'h3, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h3, 4'hf, 4'h4, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h5, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'h3, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'hf, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hd, 4'h4, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h5, 4'h4, 4'h3, 4'hf, 4'hf, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0 };
assign dw_0[107] = dw_0_107[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_108 = { 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h0, 4'h4, 4'h3, 4'h0, 4'hd, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3, 4'h3, 4'h1, 4'h5, 4'h0, 4'h4, 4'h5, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5, 4'h1, 4'h5, 4'h4, 4'h5, 4'h4, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'hf, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h5, 4'h4, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'hc, 4'hf, 4'h5, 4'h5, 4'h0, 4'h1, 4'h5, 4'h0, 4'h1, 4'h1, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h3, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h3, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h7, 4'hc, 4'h0, 4'h4, 4'h3, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h4, 4'h0, 4'h5, 4'h5, 4'h1, 4'h1, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf };
assign dw_0[108] = dw_0_108[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_109 = { 4'hc, 4'hf, 4'hc, 4'h3, 4'h0, 4'hc, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'h1, 4'h1, 4'h0, 4'h1, 4'h1, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h1, 4'h4, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'hc, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'hf, 4'hc, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h3, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h3, 4'hf, 4'h3, 4'hc, 4'h3, 4'h3, 4'hc, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h3, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h5, 4'h5, 4'h1, 4'h1, 4'h0, 4'h0, 4'h5, 4'hc, 4'h3, 4'hf, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h3, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h3, 4'hc, 4'hc, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h3, 4'hf, 4'h4, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h4, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf };
assign dw_0[109] = dw_0_109[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_110 = { 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'hf, 4'h4, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'h1, 4'h1, 4'h4, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc, 4'hc, 4'h5, 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'hc, 4'hc, 4'hc, 4'h0, 4'hc, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h5, 4'h3, 4'h1, 4'h5, 4'h3, 4'h3, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h1, 4'h1, 4'h4, 4'h3, 4'h1, 4'hc, 4'h0, 4'h1, 4'h5, 4'h4, 4'h0, 4'h1, 4'h7, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'h3, 4'hc, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'hc, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'hc, 4'h4, 4'h1, 4'h4, 4'h5, 4'h5, 4'h1, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hd, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'h0, 4'hd, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h3, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h1, 4'h3, 4'h1, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h3, 4'h4, 4'hc, 4'h3, 4'h0, 4'hc, 4'hc, 4'hf, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'hc, 4'hf, 4'hc, 4'hc, 4'h3, 4'hd, 4'h1, 4'h5, 4'h1, 4'h5, 4'h4, 4'h1, 4'h0, 4'h1, 4'hf, 4'hc, 4'h3, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h7, 4'hc, 4'h0, 4'h3, 4'hf, 4'h0, 4'h3, 4'hd };
assign dw_0[110] = dw_0_110[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_111 = { 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'hc, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'hf, 4'hc, 4'h1, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'hd, 4'h4, 4'hc, 4'h3, 4'h1, 4'h3, 4'hf, 4'h3, 4'h1, 4'h4, 4'hc, 4'h4, 4'h5, 4'h4, 4'h1, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'hf, 4'hd, 4'hc, 4'h0, 4'h0, 4'h4, 4'h5, 4'h4, 4'h0, 4'hf, 4'hd, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h1, 4'hf, 4'h5, 4'hc, 4'hc, 4'h0, 4'h0, 4'h4, 4'hc, 4'hf, 4'hc, 4'h4, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h7, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h3, 4'h5, 4'h4, 4'h1, 4'h4, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'hd, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hd, 4'h4, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h7, 4'h1, 4'h0, 4'h3, 4'h1, 4'h0, 4'hf, 4'h0, 4'h1, 4'hf, 4'h4, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'hf, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h1, 4'h1, 4'h5, 4'h3, 4'h0, 4'h7, 4'hc, 4'h3, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h3, 4'hf, 4'h0, 4'h1, 4'h0, 4'h4, 4'h4, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hd, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'hf, 4'h5, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hd, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hc, 4'hf, 4'hd, 4'hc, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd };
assign dw_0[111] = dw_0_111[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_112 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h1, 4'h4, 4'hf, 4'h1, 4'h0, 4'h3, 4'h0, 4'h4, 4'hc, 4'h3, 4'hf, 4'h0, 4'h1, 4'h1, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h5, 4'h4, 4'h1, 4'h5, 4'hf, 4'h4, 4'h0, 4'h3, 4'h7, 4'h5, 4'h4, 4'h3, 4'h0, 4'hf, 4'h1, 4'h0, 4'h1, 4'h4, 4'h4, 4'h5, 4'h1, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h1, 4'h5, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'h3, 4'h3, 4'hc, 4'hf, 4'h0, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h4, 4'h1, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h1, 4'h4, 4'hc, 4'h0, 4'h1, 4'h4, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'hc, 4'h0, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h3, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h5, 4'h0, 4'h4, 4'h0, 4'hc, 4'hc, 4'hf, 4'hc, 4'h0, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h3, 4'h0, 4'hf, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'h5, 4'h0, 4'h3, 4'h0, 4'h5, 4'h1, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h3, 4'h5, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'hc, 4'hf, 4'hf, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'hf, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3 };
assign dw_0[112] = dw_0_112[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_113 = { 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h0, 4'hc, 4'hc, 4'h1, 4'hf, 4'hc, 4'hc, 4'h3, 4'h3, 4'h0, 4'h4, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h4, 4'hf, 4'hc, 4'h0, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'h7, 4'hf, 4'h0, 4'hf, 4'hc, 4'h7, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h4, 4'hc, 4'h7, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'hf, 4'hc, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h3, 4'h0, 4'h5, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h5, 4'hf, 4'hf, 4'h3, 4'h3, 4'h3, 4'hf, 4'hc, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'h3, 4'h3, 4'h3, 4'hc, 4'hf, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h1, 4'h1, 4'h3, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'hc, 4'hf, 4'h3, 4'hf, 4'hc, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h1, 4'h1, 4'h5, 4'h1, 4'h4, 4'h5, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'h1, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h5, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'hc, 4'hc, 4'hf, 4'h3, 4'h4, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h4, 4'h1, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'hf, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h1, 4'hc, 4'hc, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'hc, 4'h4, 4'hc, 4'h1, 4'h3, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'hd, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h3 };
assign dw_0[113] = dw_0_113[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_114 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h4, 4'h1, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h5, 4'h1, 4'h4, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h3, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7, 4'hf, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h0, 4'h5, 4'h1, 4'h1, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h4, 4'h5, 4'h5, 4'h1, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h5, 4'h0, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'h4, 4'h1, 4'h5, 4'h5, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'hf, 4'h3, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'h1, 4'h4, 4'h4, 4'h5, 4'h4, 4'h5, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'hc, 4'h4, 4'h0, 4'hc, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h1, 4'h1, 4'h1, 4'h4, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h5, 4'h0, 4'h0, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h3, 4'h3, 4'h3, 4'h5, 4'h4, 4'h4, 4'h4, 4'h5, 4'h1, 4'h5, 4'h5 };
assign dw_0[114] = dw_0_114[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_115 = { 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'h4, 4'hd, 4'h4, 4'h0, 4'h4, 4'h1, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h5, 4'h1, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h4, 4'hd, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h4, 4'h5, 4'h3, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h1, 4'h0, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h1, 4'hd, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h4, 4'h3, 4'h0, 4'h3, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'h3, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h4, 4'h0, 4'h7, 4'h1, 4'h1, 4'h4, 4'h5, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h3, 4'hc, 4'h3, 4'h3, 4'h3, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'hc, 4'hc, 4'h3, 4'hc, 4'h3, 4'h3, 4'h3, 4'hc, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'h3, 4'h3, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h5, 4'h1, 4'h3, 4'h3, 4'h5, 4'hc, 4'h7, 4'h0, 4'h7, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h0, 4'h0, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'hc, 4'hf, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'hc, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h1, 4'h3, 4'h3, 4'hf, 4'hc, 4'hd, 4'hc, 4'h3, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'hc, 4'h3, 4'hf, 4'hc, 4'h3, 4'hc, 4'hf, 4'h0, 4'hc, 4'h4, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5 };
assign dw_0[115] = dw_0_115[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_116 = { 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hd, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'hf, 4'h3, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'hc, 4'h4, 4'hf, 4'h0, 4'h1, 4'h4, 4'h0, 4'h5, 4'h1, 4'h0, 4'h4, 4'h3, 4'h0, 4'hf, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h4, 4'h5, 4'h5, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h0, 4'h1, 4'h5, 4'h0, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hf, 4'h3, 4'hf, 4'hf, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h1, 4'h5, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'h0, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h4, 4'h5, 4'h4, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'hc, 4'h1, 4'h1, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h4, 4'h1, 4'h1, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'hf, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'hc, 4'hf, 4'h3, 4'h3, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'h5, 4'h5, 4'h0, 4'h5, 4'h1, 4'h5, 4'h4, 4'h5, 4'h4, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h3, 4'hc, 4'h4, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h5, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'hf, 4'hf, 4'hc, 4'hc, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h3, 4'h1, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'hc, 4'h3, 4'h0, 4'h3, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'hc, 4'h5, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h1, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h7, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'hf, 4'hc, 4'hf, 4'hc, 4'h0, 4'h3, 4'hc, 4'hc };
assign dw_0[116] = dw_0_116[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_117 = { 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'h3, 4'h0, 4'h5, 4'h5, 4'h1, 4'h5, 4'h4, 4'h1, 4'h5, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h3, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h3, 4'h1, 4'h4, 4'h4, 4'h5, 4'h0, 4'h1, 4'h4, 4'h1, 4'h4, 4'h4, 4'h4, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h5, 4'h0, 4'h5, 4'h4, 4'h1, 4'h5, 4'h0, 4'h3, 4'hc, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h5, 4'h5, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'h4, 4'h0, 4'h1, 4'hc, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h4, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'hc, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h1, 4'h0, 4'h5, 4'h0, 4'h5, 4'h1, 4'h4, 4'h0, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hc, 4'h3, 4'hc, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'hf, 4'h4, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hc, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'h4, 4'h1, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hc, 4'hf, 4'hc, 4'h3, 4'h1, 4'h0, 4'h3, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h4, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5 };
assign dw_0[117] = dw_0_117[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_118 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[118] = dw_0_118[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_119 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[119] = dw_0_119[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_120 = { 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'hc, 4'h0, 4'h1, 4'h5, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h0, 4'h4, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h5, 4'h4, 4'h4, 4'h1, 4'h1, 4'h0, 4'h4, 4'h4, 4'h7, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hc, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h4, 4'h5, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h4, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h3, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h1, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'h3, 4'hf, 4'h3, 4'h0, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h3, 4'h0, 4'hf, 4'h3, 4'hc, 4'hc, 4'hc, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h1, 4'h3, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'hc, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'hc, 4'hc, 4'hc, 4'hc, 4'hf, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h7, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h3, 4'hc, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'hc, 4'hf, 4'hc, 4'h0, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h5, 4'h5, 4'h0, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h3, 4'hc, 4'hf, 4'hf, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hc, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h3, 4'hc, 4'hc, 4'hc, 4'h4, 4'h4, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h5, 4'h0, 4'h0, 4'h3, 4'hc, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'hf, 4'h0, 4'h5, 4'h0, 4'h1, 4'h5, 4'h5, 4'h0, 4'h0 };
assign dw_0[120] = dw_0_120[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_121 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[121] = dw_0_121[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_122 = { 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[122] = dw_0_122[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_123 = { 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'h4, 4'h5, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h0, 4'hc, 4'hf, 4'hc, 4'h1, 4'h5, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'hf, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h3, 4'h3, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'h0, 4'h1, 4'h5, 4'h5, 4'h1, 4'h4, 4'h5, 4'h4, 4'h5, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'hc, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'h3, 4'hf, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'hc, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'hc, 4'h0, 4'h0, 4'hc, 4'hf, 4'hf, 4'h0, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'h4, 4'h1, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'hc, 4'hf, 4'h3, 4'h0, 4'hf, 4'hf, 4'h0, 4'hc, 4'hf, 4'h0, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hf, 4'h4, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'h0, 4'h3, 4'hc, 4'h0, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h0, 4'hc, 4'h1, 4'h0, 4'h4, 4'h5, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'hc, 4'h3, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h1, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h1, 4'h1, 4'h1, 4'h5, 4'h0, 4'h4, 4'h0, 4'h1, 4'h4, 4'h1, 4'h1, 4'h1, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0 };
assign dw_0[123] = dw_0_123[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_124 = { 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'h0, 4'h1, 4'hc, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'hc, 4'hc, 4'hf, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'hd, 4'h1, 4'h0, 4'h1, 4'h5, 4'h5, 4'h5, 4'h0, 4'h4, 4'h0, 4'h4, 4'h1, 4'h1, 4'h4, 4'hf, 4'h3, 4'h3, 4'hc, 4'hc, 4'h0, 4'hc, 4'hf, 4'h1, 4'h4, 4'h3, 4'h1, 4'h1, 4'h0, 4'h0, 4'h1, 4'hf, 4'h1, 4'h4, 4'h3, 4'h3, 4'h0, 4'h4, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'h4, 4'h0, 4'h4, 4'h0, 4'hd, 4'h1, 4'h1, 4'h3, 4'hf, 4'h3, 4'hc, 4'h3, 4'h0, 4'hf, 4'h3, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'hc, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'h1, 4'h1, 4'h1, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h5, 4'h4, 4'h1, 4'h4, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'h1, 4'hc, 4'h4, 4'h5, 4'h4, 4'h1, 4'h5, 4'h4, 4'h0, 4'h0, 4'h1, 4'h4, 4'h5, 4'h1, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h4, 4'hd, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hf, 4'hf, 4'hc, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h1, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'hf, 4'hc, 4'h0, 4'hc, 4'h3, 4'h0, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h5, 4'h0, 4'h1, 4'h5, 4'h0, 4'h5, 4'h1, 4'h5, 4'h3, 4'h3, 4'hf, 4'hf, 4'hc, 4'hf, 4'h3, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h0, 4'h5, 4'hc, 4'h5, 4'h1, 4'h0, 4'h0, 4'h4, 4'h5, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h1, 4'h4, 4'h5, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h0, 4'hf, 4'hc, 4'hc, 4'hc, 4'hc, 4'h3, 4'hc, 4'hf, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h4, 4'h0, 4'h0, 4'hf, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h3, 4'h4, 4'h3, 4'h4, 4'hf, 4'h1, 4'h5, 4'hc, 4'h4, 4'h0, 4'h4, 4'hf, 4'hf, 4'hc, 4'hc, 4'h3, 4'h0, 4'hc, 4'h3, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'h3, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h5, 4'h1, 4'h7, 4'h4, 4'h5, 4'hc, 4'h0, 4'hc, 4'h7, 4'h4, 4'h3, 4'h5, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h5, 4'h0, 4'hf, 4'hf, 4'h1, 4'h1, 4'h3, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h3, 4'h1, 4'h0, 4'h4, 4'h5, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h7 };
assign dw_0[124] = dw_0_124[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_125 = { 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h4, 4'h1, 4'h4, 4'hc, 4'h3, 4'h0, 4'h0, 4'hf, 4'hf, 4'h3, 4'h3, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'h5, 4'h4, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'h0, 4'hc, 4'hf, 4'h3, 4'h0, 4'h5, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h4, 4'h4, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'h0, 4'h5, 4'hc, 4'h3, 4'h0, 4'h0, 4'h4, 4'h4, 4'h3, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'h3, 4'h3, 4'h3, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'h3, 4'h0, 4'h3, 4'h0, 4'hf, 4'h3, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'h4, 4'h0, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h5, 4'h4, 4'h5, 4'h5, 4'h3, 4'h5, 4'h0, 4'h1, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'hf, 4'h3, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hf, 4'hc, 4'hc, 4'h0, 4'hc, 4'h3, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'h5, 4'h1, 4'h4, 4'h0, 4'h1, 4'h1, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h1, 4'h5, 4'h5, 4'h1, 4'h5, 4'hc, 4'h0, 4'h0, 4'h3, 4'hc, 4'h7, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'h1, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h7, 4'h3, 4'h3, 4'h3, 4'h0, 4'h3, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h0, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'hc, 4'hc, 4'h3, 4'hc, 4'hf, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'hd, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h1, 4'h0, 4'h3, 4'h0, 4'h1, 4'h4, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h5, 4'h4, 4'h0, 4'h1, 4'h1, 4'h1, 4'h0, 4'h4, 4'h1, 4'h1, 4'h4, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'hc, 4'hf, 4'h0, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'hf, 4'hc, 4'h0, 4'hf, 4'h3, 4'hc, 4'h4, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h0, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hf, 4'hf, 4'h0, 4'h0, 4'h4, 4'h1, 4'hd, 4'h5, 4'h3, 4'hc, 4'h0, 4'h0, 4'hf, 4'hc, 4'hc, 4'hf, 4'hc, 4'hf, 4'hc, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h3, 4'hf, 4'h0, 4'hf, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h1, 4'h1, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h4, 4'h4, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'h4, 4'h1, 4'h5, 4'h0, 4'h0, 4'h1, 4'h1, 4'h4 };
assign dw_0[125] = dw_0_125[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_126 = { 4'h0, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h4, 4'hf, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'h3, 4'h3, 4'h5, 4'h1, 4'h0, 4'h4, 4'h5, 4'h5, 4'h1, 4'h5, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h4, 4'h1, 4'h1, 4'h0, 4'h1, 4'h0, 4'hf, 4'h3, 4'hf, 4'h3, 4'h3, 4'hf, 4'hf, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h4, 4'h4, 4'h5, 4'h4, 4'h5, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h1, 4'h1, 4'h4, 4'h0, 4'h5, 4'h0, 4'h5, 4'h5, 4'h1, 4'h0, 4'h0, 4'h3, 4'hd, 4'h0, 4'h3, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'hc, 4'hf, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h4, 4'hc, 4'h3, 4'h0, 4'hf, 4'h3, 4'h3, 4'hc, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h1, 4'h5, 4'hc, 4'h0, 4'h0, 4'h0, 4'h4, 4'hc, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h1, 4'h4, 4'h1, 4'h0, 4'h0, 4'h5, 4'h1, 4'h5, 4'h4, 4'h1, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h4, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h3, 4'hf, 4'hc, 4'h0, 4'h3, 4'hf, 4'hc, 4'h0, 4'h3, 4'hc, 4'h4, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'hc, 4'h0, 4'hf, 4'hf, 4'hc, 4'h0, 4'h3, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h1, 4'h4, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h4, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h4, 4'h4, 4'h0, 4'h1, 4'h4, 4'h0, 4'h1, 4'h0, 4'h1, 4'h5, 4'h4, 4'h5, 4'h5, 4'h5, 4'h4, 4'h4, 4'h5, 4'h0, 4'h1, 4'h1, 4'h0, 4'h4, 4'h4, 4'h1, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'h0, 4'h1, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h1, 4'h1, 4'h4, 4'h1, 4'h4, 4'h4, 4'h0, 4'h5, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'hc, 4'h0, 4'h3, 4'h3, 4'hc, 4'h3, 4'hc, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h7, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hd, 4'hc, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'hc, 4'hf, 4'hf, 4'hf, 4'h0, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h1, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h5, 4'h0, 4'h4, 4'h4, 4'h5, 4'h4, 4'h4, 4'h1, 4'h4, 4'h0, 4'h1, 4'hf, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'hc };
assign dw_0[126] = dw_0_126[d0_cntr];
reg [D0_CYC-1:0][D0_IN_SIZE*D0_BW_W-1:0] dw_0_127 = { 4'hf, 4'hf, 4'h3, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h5, 4'h1, 4'h4, 4'h5, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'hc, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h4, 4'h0, 4'h4, 4'h5, 4'h5, 4'h5, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'hc, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'hf, 4'hf, 4'hf, 4'hc, 4'h3, 4'hc, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'hf, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h3, 4'h3, 4'h0, 4'hc, 4'hc, 4'hc, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'hc, 4'h3, 4'h0, 4'hf, 4'h0, 4'h3, 4'hf, 4'hc, 4'hc, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'hf, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h1, 4'h5, 4'h0, 4'h1, 4'h0, 4'h4, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'hf, 4'h0, 4'h3, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h5, 4'h4, 4'h4, 4'h0, 4'h0, 4'h5, 4'h4, 4'h0, 4'h0, 4'h0, 4'h3, 4'hf, 4'h3, 4'hc, 4'hc, 4'hf, 4'hf, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'hc, 4'h3, 4'h3, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'hc, 4'h0, 4'hc, 4'h0, 4'h0, 4'h0, 4'h0, 4'h3, 4'h0, 4'h0, 4'h0, 4'h5, 4'h1, 4'h4, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h1, 4'h5, 4'h5, 4'h5, 4'h5, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h4, 4'h5, 4'h4, 4'h5, 4'h1, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h5, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h4, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h1, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0, 4'h0 };
assign dw_0[127] = dw_0_127[d0_cntr];
