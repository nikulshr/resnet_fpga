module convlyr1 (
input clock,
input reset,
input vld_in,
input [5:0][15:0] in,
output vld_out,
output [63:0][15:0] out
);
reg [3:0] vld_reg = 0;
wire [3:0] resets;
reg [2:0] rst_reg;
assign resets = { rst_reg, reset };
assign vld_out = vld_reg[3];
always @( posedge clock ) begin
vld_reg <= { vld_reg[2:0], vld_in };
rst_reg <= resets[2:0];
end
reg [15:0] tree_0;
always @( posedge clock ) begin
tree_0 <= ( $signed( in[0] ) ) + ( $signed( in[2] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1;
always @( posedge clock ) begin
tree_1 <= ( $signed( in[4] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2;
always @( posedge clock ) begin
tree_2 <= ( $signed( tree_0 ) ) + ( $signed( tree_1 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3;
always @( posedge clock ) begin
tree_3 <= ( $signed( in[0] ) ) + ( $signed( in[2] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_4;
always @( posedge clock ) begin
tree_4 <= ( $signed( in[4] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_5;
always @( posedge clock ) begin
tree_5 <= ( $signed( tree_3 ) ) + ( $signed( tree_4 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_6;
always @( posedge clock ) begin
tree_6 <= ( $signed( in[0] ) ) - ( $signed( in[4] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_7;
always @( posedge clock ) begin
tree_7 <= ( $signed( in[2] ) ) + ( $signed( in[4] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_8;
always @( posedge clock ) begin
tree_8 <= ( $signed( in[5] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_9;
always @( posedge clock ) begin
tree_9 <= ( $signed( tree_7 ) ) + ( $signed( tree_8 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_10;
always @( posedge clock ) begin
tree_10 <= ( $signed( in[1] ) ) - ( $signed( in[5] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_11;
always @( posedge clock ) begin
tree_11 <= ( $signed( in[3] ) ) - ( $signed( in[4] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_12;
always @( posedge clock ) begin
tree_12 <= ( $signed( in[0] ) ) + ( $signed( in[2] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_13;
always @( posedge clock ) begin
tree_13 <= ( $signed( tree_6 ) ) + ( $signed( tree_10 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_14;
always @( posedge clock ) begin
tree_14 <= ( $signed( in[0] ) ) + ( $signed( in[2] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_15;
always @( posedge clock ) begin
tree_15 <= ( $signed( in[3] ) ) + ( $signed( in[4] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_16;
always @( posedge clock ) begin
tree_16 <= ( $signed( in[5] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_17;
always @( posedge clock ) begin
tree_17 <= ( $signed( tree_15 ) ) + ( $signed( tree_16 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_18;
always @( posedge clock ) begin
tree_18 <= ( $signed( in[5] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_19;
always @( posedge clock ) begin
tree_19 <= ( $signed( tree_18 ) ) + ( $signed( tree_6 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_20;
always @( posedge clock ) begin
tree_20 <= ( $signed( in[1] ) ) + ( $signed( in[3] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_21;
always @( posedge clock ) begin
tree_21 <= ( $signed( in[5] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_22;
always @( posedge clock ) begin
tree_22 <= ( $signed( tree_21 ) ) + ( $signed( tree_6 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_23;
always @( posedge clock ) begin
tree_23 <= ( $signed( tree_6 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_24;
always @( posedge clock ) begin
tree_24 <= ( $signed( tree_10 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_25;
always @( posedge clock ) begin
tree_25 <= ( $signed( in[4] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_26;
always @( posedge clock ) begin
tree_26 <= ( $signed( tree_25 ) ) - ( $signed( tree_10 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_27;
always @( posedge clock ) begin
tree_27 <= ( $signed( in[0] ) ) + ( $signed( in[2] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_28;
always @( posedge clock ) begin
tree_28 <= ( $signed( tree_27 ) ) + ( $signed( tree_10 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_29;
always @( posedge clock ) begin
tree_29 <= ( $signed( in[1] ) ) + ( $signed( in[3] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_30;
always @( posedge clock ) begin
tree_30 <= ( $signed( in[5] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_31;
always @( posedge clock ) begin
tree_31 <= ( $signed( tree_29 ) ) + ( $signed( tree_30 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_32;
always @( posedge clock ) begin
tree_32 <= ( $signed( in[0] ) ) + ( $signed( in[4] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_33;
always @( posedge clock ) begin
tree_33 <= ( $signed( in[1] ) ) + ( $signed( in[3] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_34;
always @( posedge clock ) begin
tree_34 <= ( $signed( in[1] ) ) - ( $signed( in[2] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_35;
always @( posedge clock ) begin
tree_35 <= ( $signed( in[5] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_36;
always @( posedge clock ) begin
tree_36 <= ( $signed( tree_35 ) ) + ( $signed( tree_6 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_37;
always @( posedge clock ) begin
tree_37 <= ( $signed( in[3] ) ) + ( $signed( in[5] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_38;
always @( posedge clock ) begin
tree_38 <= ( $signed( in[1] ) ) + ( $signed( in[3] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_39;
always @( posedge clock ) begin
tree_39 <= ( $signed( tree_6 ) ) + ( $signed( tree_10 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_40;
always @( posedge clock ) begin
tree_40 <= ( $signed( in[0] ) ) + ( $signed( in[1] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_41;
always @( posedge clock ) begin
tree_41 <= ( $signed( in[2] ) ) + ( $signed( in[3] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_42;
always @( posedge clock ) begin
tree_42 <= ( $signed( tree_40 ) ) + ( $signed( tree_41 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_43;
always @( posedge clock ) begin
tree_43 <= ( $signed( tree_34 ) ) - ( $signed( tree_11 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_44;
always @( posedge clock ) begin
tree_44 <= ( $signed( in[1] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_45;
always @( posedge clock ) begin
tree_45 <= ( $signed( in[0] ) ) + ( $signed( in[2] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_46;
always @( posedge clock ) begin
tree_46 <= ( $signed( in[4] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_47;
always @( posedge clock ) begin
tree_47 <= ( $signed( tree_45 ) ) + ( $signed( tree_46 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_48;
always @( posedge clock ) begin
tree_48 <= ( $signed( in[1] ) ) + ( $signed( in[3] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_49;
always @( posedge clock ) begin
tree_49 <= ( $signed( in[1] ) ) + ( $signed( in[2] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_50;
always @( posedge clock ) begin
tree_50 <= ( $signed( in[3] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_51;
always @( posedge clock ) begin
tree_51 <= ( $signed( tree_49 ) ) + ( $signed( tree_50 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_52;
always @( posedge clock ) begin
tree_52 <= ( $signed( in[4] ) ) - ( $signed( in[5] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_53;
always @( posedge clock ) begin
tree_53 <= ( $signed( in[5] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_54;
always @( posedge clock ) begin
tree_54 <= ( $signed( tree_6 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_55;
always @( posedge clock ) begin
tree_55 <= ( $signed( in[1] ) ) + ( $signed( in[3] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_56;
always @( posedge clock ) begin
tree_56 <= ( $signed( in[5] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_57;
always @( posedge clock ) begin
tree_57 <= ( $signed( in[0] ) ) - ( $signed( in[5] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_58;
always @( posedge clock ) begin
tree_58 <= ( $signed( in[3] ) ) + ( $signed( in[5] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_59;
always @( posedge clock ) begin
tree_59 <= ( $signed( in[0] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_60;
always @( posedge clock ) begin
tree_60 <= ( $signed( tree_59 ) ) - ( $signed( tree_10 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_61;
always @( posedge clock ) begin
tree_61 <= ( $signed( in[0] ) ) + ( $signed( in[2] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_62;
always @( posedge clock ) begin
tree_62 <=  - ( $signed( tree_61 ) ) + ( $signed( tree_11 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_63;
always @( posedge clock ) begin
tree_63 <= ( $signed( in[0] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_64;
always @( posedge clock ) begin
tree_64 <= ( $signed( in[0] ) ) - ( $signed( in[3] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_65;
always @( posedge clock ) begin
tree_65 <= ( $signed( tree_64 ) ) - ( $signed( tree_34 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_66;
always @( posedge clock ) begin
tree_66 <= ( $signed( in[1] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_67;
always @( posedge clock ) begin
tree_67 <= ( $signed( in[0] ) ) + ( $signed( in[2] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_68;
always @( posedge clock ) begin
tree_68 <= ( $signed( in[0] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_69;
always @( posedge clock ) begin
tree_69 <= ( $signed( tree_10 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_70;
always @( posedge clock ) begin
tree_70 <= ( $signed( in[4] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_71;
always @( posedge clock ) begin
tree_71 <= ( $signed( in[1] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_72;
always @( posedge clock ) begin
tree_72 <= ( $signed( in[1] ) ) + ( $signed( in[5] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_73;
always @( posedge clock ) begin
tree_73 <= ( $signed( in[1] ) ) + ( $signed( in[3] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_74;
always @( posedge clock ) begin
tree_74 <= ( $signed( in[5] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_75;
always @( posedge clock ) begin
tree_75 <= ( $signed( tree_73 ) ) + ( $signed( tree_74 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_76;
always @( posedge clock ) begin
tree_76 <= ( $signed( in[2] ) ) + ( $signed( in[4] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_77;
always @( posedge clock ) begin
tree_77 <= ( $signed( in[2] ) ) + ( $signed( in[4] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_78;
always @( posedge clock ) begin
tree_78 <= ( $signed( tree_26 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_79;
always @( posedge clock ) begin
tree_79 <= ( $signed( in[0] ) ) + ( $signed( in[2] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_80;
always @( posedge clock ) begin
tree_80 <= ( $signed( in[1] ) ) + ( $signed( in[3] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_81;
always @( posedge clock ) begin
tree_81 <= ( $signed( tree_52 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_82;
always @( posedge clock ) begin
tree_82 <= ( $signed( in[0] ) ) + ( $signed( in[2] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_83;
always @( posedge clock ) begin
tree_83 <= ( $signed( tree_57 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_84;
always @( posedge clock ) begin
tree_84 <= ( $signed( in[0] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_85;
always @( posedge clock ) begin
tree_85 <= ( $signed( in[5] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_86;
always @( posedge clock ) begin
tree_86 <= ( $signed( tree_85 ) ) - ( $signed( tree_6 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_87;
always @( posedge clock ) begin
tree_87 <= ( $signed( tree_6 ) ) - ( $signed( tree_10 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_88;
always @( posedge clock ) begin
tree_88 <= ( $signed( in[1] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_89;
always @( posedge clock ) begin
tree_89 <= ( $signed( tree_88 ) ) + ( $signed( tree_11 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_90;
always @( posedge clock ) begin
tree_90 <= ( $signed( in[3] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_91;
always @( posedge clock ) begin
tree_91 <= ( $signed( tree_90 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_92;
always @( posedge clock ) begin
tree_92 <= ( $signed( tree_91 ) ) + ( $signed( tree_86 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_93;
always @( posedge clock ) begin
tree_93 <= ( $signed( tree_26 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_94;
always @( posedge clock ) begin
tree_94 <= ( $signed( in[3] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_95;
always @( posedge clock ) begin
tree_95 <= ( $signed( tree_94 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_96;
always @( posedge clock ) begin
tree_96 <= ( $signed( tree_95 ) ) + ( $signed( tree_86 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_97;
always @( posedge clock ) begin
tree_97 <= ( $signed( in[4] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_98;
always @( posedge clock ) begin
tree_98 <= ( $signed( tree_97 ) ) - ( $signed( tree_34 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_99;
always @( posedge clock ) begin
tree_99 <= ( $signed( tree_87 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_100;
always @( posedge clock ) begin
tree_100 <= ( $signed( in[2] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_101;
always @( posedge clock ) begin
tree_101 <= ( $signed( tree_100 ) ) + ( $signed( tree_52 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_102;
always @( posedge clock ) begin
tree_102 <= ( $signed( tree_87 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_103;
always @( posedge clock ) begin
tree_103 <= ( $signed( in[2] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_104;
always @( posedge clock ) begin
tree_104 <= ( $signed( tree_103 ) ) + ( $signed( tree_57 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_105;
always @( posedge clock ) begin
tree_105 <= ( $signed( tree_86 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_106;
always @( posedge clock ) begin
tree_106 <= ( $signed( tree_87 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_107;
always @( posedge clock ) begin
tree_107 <=  - ( $signed( tree_9 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_108;
always @( posedge clock ) begin
tree_108 <=  - ( $signed( tree_13 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_109;
always @( posedge clock ) begin
tree_109 <=  - ( $signed( tree_14 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_110;
always @( posedge clock ) begin
tree_110 <=  - ( $signed( tree_22 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_111;
always @( posedge clock ) begin
tree_111 <=  - ( $signed( tree_24 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_112;
always @( posedge clock ) begin
tree_112 <=  - ( $signed( tree_28 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_113;
always @( posedge clock ) begin
tree_113 <=  - ( $signed( tree_31 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_114;
always @( posedge clock ) begin
tree_114 <=  - ( $signed( tree_33 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_115;
always @( posedge clock ) begin
tree_115 <=  - ( $signed( tree_36 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_116;
always @( posedge clock ) begin
tree_116 <=  - ( $signed( tree_37 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_117;
always @( posedge clock ) begin
tree_117 <=  - ( $signed( tree_38 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_118;
always @( posedge clock ) begin
tree_118 <=  - ( $signed( tree_42 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_119;
always @( posedge clock ) begin
tree_119 <=  - ( $signed( tree_47 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_120;
always @( posedge clock ) begin
tree_120 <=  - ( $signed( tree_48 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_121;
always @( posedge clock ) begin
tree_121 <=  - ( $signed( tree_54 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_122;
always @( posedge clock ) begin
tree_122 <=  - ( $signed( tree_55 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_123;
always @( posedge clock ) begin
tree_123 <=  - ( $signed( tree_58 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_124;
always @( posedge clock ) begin
tree_124 <=  - ( $signed( tree_68 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_125;
always @( posedge clock ) begin
tree_125 <=  - ( $signed( tree_70 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_126;
always @( posedge clock ) begin
tree_126 <=  - ( $signed( tree_71 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_127;
always @( posedge clock ) begin
tree_127 <=  - ( $signed( tree_76 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_128;
always @( posedge clock ) begin
tree_128 <=  - ( $signed( tree_77 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_129;
always @( posedge clock ) begin
tree_129 <=  - ( $signed( tree_78 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_130;
always @( posedge clock ) begin
tree_130 <=  - ( $signed( tree_80 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_131;
always @( posedge clock ) begin
tree_131 <=  - ( $signed( tree_81 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_132;
always @( posedge clock ) begin
tree_132 <=  - ( $signed( tree_82 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_133;
always @( posedge clock ) begin
tree_133 <=  - ( $signed( tree_83 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_134;
always @( posedge clock ) begin
tree_134 <=  - ( $signed( tree_92 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_135;
always @( posedge clock ) begin
tree_135 <=  - ( $signed( tree_99 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_136;
always @( posedge clock ) begin
tree_136 <=  - ( $signed( tree_105 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_137;
always @( posedge clock ) begin
tree_137 <=  - ( $signed( tree_106 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [1:0][15:0] out_0;
assign out[0] = out_0[1];
reg [1:0][15:0] out_1;
assign out[1] = out_1[1];
assign out[2] = tree_136;
reg [15:0] out_3;
assign out[3] = out_3;
assign out[4] = tree_137;
reg [1:0][15:0] out_5;
assign out[5] = out_5[1];
reg [2:0][15:0] out_6;
assign out[6] = out_6[2];
reg [15:0] out_7;
assign out[7] = out_7;
assign out[8] = tree_134;
reg [1:0][15:0] out_9;
assign out[9] = out_9[1];
reg [1:0][15:0] out_10;
assign out[10] = out_10[1];
reg [1:0][15:0] out_11;
assign out[11] = out_11[1];
reg [2:0][15:0] out_12;
assign out[12] = out_12[2];
reg [15:0] out_13;
assign out[13] = out_13;
reg [1:0][15:0] out_14;
assign out[14] = out_14[1];
reg [15:0] out_15;
assign out[15] = out_15;
reg [15:0] out_16;
assign out[16] = out_16;
reg [15:0] out_17;
assign out[17] = out_17;
reg [15:0] out_18;
assign out[18] = out_18;
reg [15:0] out_19;
assign out[19] = out_19;
reg [2:0][15:0] out_20;
assign out[20] = out_20[2];
reg [1:0][15:0] out_21;
assign out[21] = out_21[1];
reg [1:0][15:0] out_22;
assign out[22] = out_22[1];
reg [15:0] out_23;
assign out[23] = out_23;
assign out[24] = tree_135;
reg [1:0][15:0] out_25;
assign out[25] = out_25[1];
reg [1:0][15:0] out_26;
assign out[26] = out_26[1];
reg [1:0][15:0] out_27;
assign out[27] = out_27[1];
reg [15:0] out_28;
assign out[28] = out_28;
reg [1:0][15:0] out_29;
assign out[29] = out_29[1];
reg [2:0][15:0] out_30;
assign out[30] = out_30[2];
reg [15:0] out_31;
assign out[31] = out_31;
reg [1:0][15:0] out_32;
assign out[32] = out_32[1];
reg [1:0][15:0] out_33;
assign out[33] = out_33[1];
reg [1:0][15:0] out_34;
assign out[34] = out_34[1];
reg [2:0][15:0] out_35;
assign out[35] = out_35[2];
reg [15:0] out_36;
assign out[36] = out_36;
reg [1:0][15:0] out_37;
assign out[37] = out_37[1];
reg [2:0][15:0] out_38;
assign out[38] = out_38[2];
reg [15:0] out_39;
assign out[39] = out_39;
reg [1:0][15:0] out_40;
assign out[40] = out_40[1];
reg [1:0][15:0] out_41;
assign out[41] = out_41[1];
reg [1:0][15:0] out_42;
assign out[42] = out_42[1];
reg [1:0][15:0] out_43;
assign out[43] = out_43[1];
reg [2:0][15:0] out_44;
assign out[44] = out_44[2];
reg [1:0][15:0] out_45;
assign out[45] = out_45[1];
reg [2:0][15:0] out_46;
assign out[46] = out_46[2];
reg [2:0][15:0] out_47;
assign out[47] = out_47[2];
reg [1:0][15:0] out_48;
assign out[48] = out_48[1];
reg [1:0][15:0] out_49;
assign out[49] = out_49[1];
reg [1:0][15:0] out_50;
assign out[50] = out_50[1];
reg [1:0][15:0] out_51;
assign out[51] = out_51[1];
reg [2:0][15:0] out_52;
assign out[52] = out_52[2];
reg [1:0][15:0] out_53;
assign out[53] = out_53[1];
reg [1:0][15:0] out_54;
assign out[54] = out_54[1];
assign out[55] = 16'h0;
reg [1:0][15:0] out_56;
assign out[56] = out_56[1];
assign out[57] = tree_129;
reg [2:0][15:0] out_58;
assign out[58] = out_58[2];
reg [1:0][15:0] out_59;
assign out[59] = out_59[1];
reg [15:0] out_60;
assign out[60] = out_60;
reg [1:0][15:0] out_61;
assign out[61] = out_61[1];
reg [15:0] out_62;
assign out[62] = out_62;
reg [2:0][15:0] out_63;
assign out[63] = out_63[2];
always @( posedge clock ) begin
out_0 <= { out_0[0:0], tree_2};
out_1 <= { out_1[0:0], tree_5};
out_3 <= tree_107;
out_5 <= { out_5[0:0], tree_89};
out_6 <= { out_6[1:0], tree_12};
out_7 <= tree_108;
out_9 <= { out_9[0:0], tree_109};
out_10 <= { out_10[0:0], tree_17};
out_11 <= { out_11[0:0], tree_19};
out_12 <= { out_12[1:0], tree_20};
out_13 <= tree_110;
out_14 <= { out_14[0:0], tree_23};
out_15 <= tree_111;
out_16 <= tree_93;
out_17 <= tree_112;
out_18 <= tree_113;
out_19 <= tree_96;
out_20 <= { out_20[1:0], tree_32};
out_21 <= { out_21[0:0], tree_114};
out_22 <= { out_22[0:0], tree_98};
out_23 <= tree_115;
out_25 <= { out_25[0:0], tree_116};
out_26 <= { out_26[0:0], tree_117};
out_27 <= { out_27[0:0], tree_39};
out_28 <= tree_118;
out_29 <= { out_29[0:0], tree_43};
out_30 <= { out_30[1:0], tree_44};
out_31 <= tree_119;
out_32 <= { out_32[0:0], tree_120};
out_33 <= { out_33[0:0], tree_51};
out_34 <= { out_34[0:0], tree_101};
out_35 <= { out_35[1:0], tree_53};
out_36 <= tree_121;
out_37 <= { out_37[0:0], tree_122};
out_38 <= { out_38[1:0], tree_56};
out_39 <= tree_102;
out_40 <= { out_40[0:0], tree_104};
out_41 <= { out_41[0:0], tree_123};
out_42 <= { out_42[0:0], tree_60};
out_43 <= { out_43[0:0], tree_62};
out_44 <= { out_44[1:0], tree_63};
out_45 <= { out_45[0:0], tree_65};
out_46 <= { out_46[1:0], tree_66};
out_47 <= { out_47[1:0], tree_67};
out_48 <= { out_48[0:0], tree_124};
out_49 <= { out_49[0:0], tree_69};
out_50 <= { out_50[0:0], tree_125};
out_51 <= { out_51[0:0], tree_126};
out_52 <= { out_52[1:0], tree_72};
out_53 <= { out_53[0:0], tree_75};
out_54 <= { out_54[0:0], tree_127};
out_56 <= { out_56[0:0], tree_128};
out_58 <= { out_58[1:0], tree_79};
out_59 <= { out_59[0:0], tree_130};
out_60 <= tree_131;
out_61 <= { out_61[0:0], tree_132};
out_62 <= tree_133;
out_63 <= { out_63[1:0], tree_84};
end
endmodule
