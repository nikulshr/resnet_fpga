localparam D2_IN_SIZE = 1;
localparam D2_BW_W = 16;
localparam D2_SHIFT = 6;
localparam LOG2_D2_CYC = 5;
localparam D2_CYC = 24;
localparam D2_CH = 128;
reg [LOG2_D2_CYC-1:0] d2_cntr;
wire [D2_CH-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2;
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_0 = { 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'h0040, 16'hffc0, 16'h0000, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0040, 16'hffc0 };
assign dw_2[0] = dw_2_0[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_1 = { 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'h0040 };
assign dw_2[1] = dw_2_1[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_2 = { 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'h0040, 16'h0040, 16'h0040, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0 };
assign dw_2[2] = dw_2_2[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_3 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[3] = dw_2_3[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_4 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[4] = dw_2_4[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_5 = { 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[5] = dw_2_5[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_6 = { 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000 };
assign dw_2[6] = dw_2_6[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_7 = { 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0 };
assign dw_2[7] = dw_2_7[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_8 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000 };
assign dw_2[8] = dw_2_8[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_9 = { 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0040, 16'h0000, 16'h0040, 16'h0000, 16'hffc0, 16'h0040 };
assign dw_2[9] = dw_2_9[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_10 = { 16'hffc0, 16'h0040, 16'h0000, 16'h0040, 16'h0040, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0 };
assign dw_2[10] = dw_2_10[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_11 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[11] = dw_2_11[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_12 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[12] = dw_2_12[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_13 = { 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000 };
assign dw_2[13] = dw_2_13[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_14 = { 16'hffc0, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000 };
assign dw_2[14] = dw_2_14[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_15 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[15] = dw_2_15[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_16 = { 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'h0040, 16'h0040 };
assign dw_2[16] = dw_2_16[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_17 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[17] = dw_2_17[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_18 = { 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'h0040, 16'h0040, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0040 };
assign dw_2[18] = dw_2_18[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_19 = { 16'h0040, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000 };
assign dw_2[19] = dw_2_19[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_20 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000 };
assign dw_2[20] = dw_2_20[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_21 = { 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'hffc0, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0 };
assign dw_2[21] = dw_2_21[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_22 = { 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0000 };
assign dw_2[22] = dw_2_22[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_23 = { 16'h0000, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[23] = dw_2_23[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_24 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[24] = dw_2_24[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_25 = { 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0040 };
assign dw_2[25] = dw_2_25[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_26 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[26] = dw_2_26[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_27 = { 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0 };
assign dw_2[27] = dw_2_27[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_28 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[28] = dw_2_28[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_29 = { 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0040 };
assign dw_2[29] = dw_2_29[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_30 = { 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[30] = dw_2_30[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_31 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[31] = dw_2_31[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_32 = { 16'h0000, 16'hffc0, 16'h0040, 16'hffc0, 16'hffc0, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0040, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'h0040 };
assign dw_2[32] = dw_2_32[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_33 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[33] = dw_2_33[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_34 = { 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[34] = dw_2_34[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_35 = { 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'hffc0, 16'h0040, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000 };
assign dw_2[35] = dw_2_35[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_36 = { 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[36] = dw_2_36[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_37 = { 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000 };
assign dw_2[37] = dw_2_37[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_38 = { 16'h0040, 16'h0000, 16'h0040, 16'h0040, 16'h0040, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000 };
assign dw_2[38] = dw_2_38[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_39 = { 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[39] = dw_2_39[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_40 = { 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0040, 16'h0040, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[40] = dw_2_40[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_41 = { 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[41] = dw_2_41[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_42 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[42] = dw_2_42[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_43 = { 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0000 };
assign dw_2[43] = dw_2_43[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_44 = { 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0040 };
assign dw_2[44] = dw_2_44[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_45 = { 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0040, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[45] = dw_2_45[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_46 = { 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000 };
assign dw_2[46] = dw_2_46[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_47 = { 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0 };
assign dw_2[47] = dw_2_47[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_48 = { 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'h0040, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[48] = dw_2_48[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_49 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0040 };
assign dw_2[49] = dw_2_49[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_50 = { 16'h0040, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0000, 16'h0040, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'hffc0, 16'hffc0, 16'h0040 };
assign dw_2[50] = dw_2_50[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_51 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[51] = dw_2_51[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_52 = { 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'hffc0, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0040, 16'hffc0, 16'hffc0 };
assign dw_2[52] = dw_2_52[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_53 = { 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0040 };
assign dw_2[53] = dw_2_53[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_54 = { 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0 };
assign dw_2[54] = dw_2_54[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_55 = { 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'hffc0, 16'hffc0, 16'h0040, 16'hffc0, 16'hffc0, 16'h0040, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000 };
assign dw_2[55] = dw_2_55[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_56 = { 16'h0040, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[56] = dw_2_56[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_57 = { 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'hffc0, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0 };
assign dw_2[57] = dw_2_57[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_58 = { 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0 };
assign dw_2[58] = dw_2_58[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_59 = { 16'h0000, 16'h0040, 16'hffc0, 16'h0040, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'h0040, 16'hffc0, 16'h0040, 16'hffc0, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000 };
assign dw_2[59] = dw_2_59[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_60 = { 16'h0040, 16'hffc0, 16'h0000, 16'h0040, 16'h0040, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'h0040, 16'h0040 };
assign dw_2[60] = dw_2_60[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_61 = { 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0040, 16'h0000 };
assign dw_2[61] = dw_2_61[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_62 = { 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0040, 16'h0000 };
assign dw_2[62] = dw_2_62[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_63 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[63] = dw_2_63[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_64 = { 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[64] = dw_2_64[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_65 = { 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0 };
assign dw_2[65] = dw_2_65[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_66 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[66] = dw_2_66[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_67 = { 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'hffc0, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0 };
assign dw_2[67] = dw_2_67[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_68 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0 };
assign dw_2[68] = dw_2_68[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_69 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[69] = dw_2_69[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_70 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0040 };
assign dw_2[70] = dw_2_70[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_71 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0000 };
assign dw_2[71] = dw_2_71[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_72 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[72] = dw_2_72[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_73 = { 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'hffc0, 16'h0000 };
assign dw_2[73] = dw_2_73[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_74 = { 16'h0040, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000 };
assign dw_2[74] = dw_2_74[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_75 = { 16'h0000, 16'h0040, 16'h0000, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000 };
assign dw_2[75] = dw_2_75[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_76 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'hffc0, 16'hffc0 };
assign dw_2[76] = dw_2_76[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_77 = { 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[77] = dw_2_77[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_78 = { 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0040 };
assign dw_2[78] = dw_2_78[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_79 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[79] = dw_2_79[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_80 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[80] = dw_2_80[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_81 = { 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000 };
assign dw_2[81] = dw_2_81[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_82 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[82] = dw_2_82[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_83 = { 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000 };
assign dw_2[83] = dw_2_83[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_84 = { 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[84] = dw_2_84[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_85 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[85] = dw_2_85[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_86 = { 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0 };
assign dw_2[86] = dw_2_86[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_87 = { 16'hffc0, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0040, 16'hffc0, 16'h0040, 16'hffc0, 16'h0040, 16'h0040, 16'hffc0, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[87] = dw_2_87[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_88 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000 };
assign dw_2[88] = dw_2_88[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_89 = { 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'hffc0, 16'hffc0, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000 };
assign dw_2[89] = dw_2_89[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_90 = { 16'hffc0, 16'hffc0, 16'hffc0, 16'h0040, 16'hffc0, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0040 };
assign dw_2[90] = dw_2_90[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_91 = { 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0000 };
assign dw_2[91] = dw_2_91[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_92 = { 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000 };
assign dw_2[92] = dw_2_92[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_93 = { 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0040 };
assign dw_2[93] = dw_2_93[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_94 = { 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0040 };
assign dw_2[94] = dw_2_94[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_95 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[95] = dw_2_95[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_96 = { 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[96] = dw_2_96[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_97 = { 16'h0000, 16'h0040, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0040 };
assign dw_2[97] = dw_2_97[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_98 = { 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[98] = dw_2_98[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_99 = { 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000 };
assign dw_2[99] = dw_2_99[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_100 = { 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'hffc0, 16'h0040 };
assign dw_2[100] = dw_2_100[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_101 = { 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[101] = dw_2_101[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_102 = { 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[102] = dw_2_102[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_103 = { 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000 };
assign dw_2[103] = dw_2_103[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_104 = { 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'h0040, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0 };
assign dw_2[104] = dw_2_104[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_105 = { 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'hffc0, 16'h0040, 16'hffc0, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0 };
assign dw_2[105] = dw_2_105[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_106 = { 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[106] = dw_2_106[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_107 = { 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0000 };
assign dw_2[107] = dw_2_107[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_108 = { 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0040 };
assign dw_2[108] = dw_2_108[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_109 = { 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'hffc0, 16'hffc0, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0 };
assign dw_2[109] = dw_2_109[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_110 = { 16'h0040, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0 };
assign dw_2[110] = dw_2_110[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_111 = { 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0040 };
assign dw_2[111] = dw_2_111[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_112 = { 16'hffc0, 16'h0040, 16'h0040, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[112] = dw_2_112[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_113 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[113] = dw_2_113[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_114 = { 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[114] = dw_2_114[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_115 = { 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0040, 16'hffc0, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[115] = dw_2_115[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_116 = { 16'hffc0, 16'h0000, 16'h0040, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0 };
assign dw_2[116] = dw_2_116[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_117 = { 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'hffc0, 16'hffc0, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[117] = dw_2_117[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_118 = { 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0040 };
assign dw_2[118] = dw_2_118[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_119 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[119] = dw_2_119[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_120 = { 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0040, 16'h0000, 16'h0040, 16'hffc0, 16'hffc0, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'h0000, 16'h0040, 16'h0040 };
assign dw_2[120] = dw_2_120[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_121 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[121] = dw_2_121[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_122 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[122] = dw_2_122[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_123 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[123] = dw_2_123[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_124 = { 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h0040, 16'h0000, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0, 16'hffc0, 16'h0000, 16'hffc0, 16'hffc0, 16'hffc0 };
assign dw_2[124] = dw_2_124[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_125 = { 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0040, 16'h0040, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[125] = dw_2_125[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_126 = { 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'hffc0, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0040, 16'h0040, 16'hffc0 };
assign dw_2[126] = dw_2_126[d2_cntr];
reg [D2_CYC-1:0][D2_IN_SIZE*D2_BW_W-1:0] dw_2_127 = { 16'h0000, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'h0000, 16'hffc0, 16'h0000, 16'h0040, 16'h0000, 16'h0000, 16'h0000, 16'h0000 };
assign dw_2[127] = dw_2_127[d2_cntr];
