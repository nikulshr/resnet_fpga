localparam BN11_CH = 64;
localparam BN11_BW_A = 4;
localparam BN11_BW_B = 15;
localparam BN11_RSHIFT = 8;
localparam BN11_BW_IN = 16;
localparam BN11_BW_OUT = 1;
localparam BN11_MAXVAL = 1;
reg [BN11_CH-1:0][BN11_BW_A-1:0] bn11_a = { 4'h3, 4'h5, 4'h5, 4'h4, 4'h4, 4'h4, 4'h6, 4'h4, 4'h4, 4'h4, 4'h5, 4'h4, 4'h6, 4'h5, 4'h5, 4'h5, 4'h4, 4'h5, 4'h5, 4'h4, 4'h4, 4'h4, 4'h4, 4'h4, 4'h4, 4'h5, 4'h4, 4'h4, 4'h4, 4'h3, 4'h3, 4'h7, 4'h5, 4'h4, 4'h4, 4'h6, 4'h3, 4'h4, 4'h5, 4'h6, 4'h5, 4'h4, 4'h6, 4'h5, 4'h4, 4'h4, 4'h5, 4'h4, 4'h4, 4'h4, 4'h4, 4'h3, 4'h4, 4'h4, 4'h4, 4'h5, 4'h4, 4'h5, 4'h6, 4'h5, 4'h4, 4'h4, 4'h4, 4'h4 };
reg [BN11_CH-1:0][BN11_BW_B-1:0] bn11_b = { 15'h6ea4, 15'h6620, 15'h7708, 15'h74a1, 15'h7687, 15'h7057, 15'h6e96, 15'h7776, 15'h74bd, 15'h7b92, 15'h717e, 15'h6fb7, 15'h62a7, 15'h683b, 15'h7a41, 15'h7f24, 15'h7036, 15'h70af, 15'h688f, 15'h752a, 15'h73a8, 15'h6cbd, 15'h6d65, 15'h718b, 15'h73f9, 15'h61bc, 15'h6ff0, 15'h76bf, 15'h7722, 15'h6a4f, 15'h7f84, 15'h5557, 15'h6dc8, 15'h76fe, 15'h7164, 15'h675f, 15'h757c, 15'h7a5d, 15'h7a3b, 15'h668a, 15'h74b6, 15'h6c65, 15'h74ec, 15'h7239, 15'h729e, 15'h7731, 15'h6ac1, 15'h6b6a, 15'h02bb, 15'h62a9, 15'h6a46, 15'h059c, 15'h6b8d, 15'h79e0, 15'h75eb, 15'h7a0b, 15'h7727, 15'h65d9, 15'h65ec, 15'h74df, 15'h6f96, 15'h6922, 15'h7958, 15'h715c };
