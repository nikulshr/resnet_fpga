localparam BN15_CH = 64;
localparam BN15_BW_A = 5;
localparam BN15_BW_B = 15;
localparam BN15_RSHIFT = 8;
localparam BN15_BW_IN = 16;
localparam BN15_BW_OUT = 1;
localparam BN15_MAXVAL = 1;
reg [BN15_CH-1:0][BN15_BW_A-1:0] bn15_a = { 5'h06, 5'h06, 5'h08, 5'h0a, 5'h06, 5'h09, 5'h05, 5'h06, 5'h08, 5'h04, 5'h0a, 5'h09, 5'h07, 5'h0a, 5'h09, 5'h09, 5'h07, 5'h05, 5'h0c, 5'h09, 5'h06, 5'h09, 5'h06, 5'h07, 5'h08, 5'h0b, 5'h08, 5'h07, 5'h08, 5'h03, 5'h06, 5'h06, 5'h0d, 5'h06, 5'h09, 5'h09, 5'h07, 5'h09, 5'h04, 5'h06, 5'h09, 5'h09, 5'h09, 5'h08, 5'h08, 5'h0b, 5'h08, 5'h08, 5'h09, 5'h07, 5'h08, 5'h0a, 5'h06, 5'h05, 5'h07, 5'h05, 5'h07, 5'h03, 5'h0a, 5'h05, 5'h09, 5'h05, 5'h06, 5'h08 };
reg [BN15_CH-1:0][BN15_BW_B-1:0] bn15_b = { 15'h0706, 15'h0a4e, 15'h0b7f, 15'h7a43, 15'h7bfb, 15'h7405, 15'h780e, 15'h7548, 15'h08f5, 15'h7f09, 15'h02b0, 15'h6b17, 15'h063e, 15'h1609, 15'h7024, 15'h310f, 15'h1c4e, 15'h7fe4, 15'h1562, 15'h4273, 15'h00e6, 15'h1149, 15'h06fc, 15'h0f2f, 15'h00eb, 15'h22b6, 15'h7bea, 15'h1106, 15'h1a78, 15'h7d1e, 15'h14e9, 15'h7e2d, 15'h0a18, 15'h2003, 15'h7e42, 15'h0d5e, 15'h0a08, 15'h7317, 15'h7fee, 15'h0c3a, 15'h7ad1, 15'h0f4e, 15'h07ee, 15'h1f8b, 15'h7955, 15'h14cc, 15'h0151, 15'h1139, 15'h71e8, 15'h0207, 15'h082b, 15'h64af, 15'h7a2d, 15'h04aa, 15'h1a06, 15'h04e4, 15'h02cb, 15'h0395, 15'h7a79, 15'h7f72, 15'h153d, 15'h05e9, 15'h7cab, 15'h77dc };
