module convlyr7 (
input clock,
input reset,
input vld_in,
input [191:0][15:0] in,
output vld_out,
output [63:0][15:0] out
);
reg [7:0] vld_reg = 0;
wire [7:0] resets;
reg [6:0] rst_reg;
assign resets = { rst_reg, reset };
assign vld_out = vld_reg[7];
always @( posedge clock ) begin
vld_reg <= { vld_reg[6:0], vld_in };
rst_reg <= resets[6:0];
end
reg [15:0] tree_0;
always @( posedge clock ) begin
tree_0 <= ( $signed( in[124] ) ) + ( $signed( in[152] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1;
always @( posedge clock ) begin
tree_1 <= ( $signed( in[161] ) ) + ( $signed( in[174] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2;
always @( posedge clock ) begin
tree_2 <= ( $signed( in[1] ) ) - ( $signed( in[21] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3;
always @( posedge clock ) begin
tree_3 <= ( $signed( in[130] ) ) - ( $signed( in[175] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_4;
always @( posedge clock ) begin
tree_4 <= ( $signed( in[87] ) ) + ( $signed( in[123] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_5;
always @( posedge clock ) begin
tree_5 <= ( $signed( in[18] ) ) + ( $signed( in[57] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_6;
always @( posedge clock ) begin
tree_6 <= ( $signed( in[22] ) ) + ( $signed( in[94] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_7;
always @( posedge clock ) begin
tree_7 <= ( $signed( in[153] ) ) + ( $signed( in[169] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_8;
always @( posedge clock ) begin
tree_8 <= ( $signed( in[72] ) ) - ( $signed( in[191] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_9;
always @( posedge clock ) begin
tree_9 <= ( $signed( in[143] ) ) - ( $signed( in[170] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_10;
always @( posedge clock ) begin
tree_10 <= ( $signed( in[43] ) ) + ( $signed( in[107] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_11;
always @( posedge clock ) begin
tree_11 <= ( $signed( in[160] ) ) + ( $signed( in[177] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_12;
always @( posedge clock ) begin
tree_12 <= ( $signed( in[112] ) ) - ( $signed( in[145] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_13;
always @( posedge clock ) begin
tree_13 <= ( $signed( in[51] ) ) + ( $signed( in[53] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_14;
always @( posedge clock ) begin
tree_14 <= ( $signed( in[120] ) ) - ( $signed( in[137] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_15;
always @( posedge clock ) begin
tree_15 <= ( $signed( in[26] ) ) - ( $signed( in[37] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_16;
always @( posedge clock ) begin
tree_16 <= ( $signed( in[7] ) ) - ( $signed( in[70] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_17;
always @( posedge clock ) begin
tree_17 <= ( $signed( in[4] ) ) + ( $signed( in[92] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_18;
always @( posedge clock ) begin
tree_18 <= ( $signed( in[90] ) ) + ( $signed( in[111] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_19;
always @( posedge clock ) begin
tree_19 <= ( $signed( in[39] ) ) - ( $signed( in[67] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_20;
always @( posedge clock ) begin
tree_20 <= ( $signed( in[133] ) ) + ( $signed( in[158] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_21;
always @( posedge clock ) begin
tree_21 <= ( $signed( in[42] ) ) + ( $signed( in[54] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_22;
always @( posedge clock ) begin
tree_22 <= ( $signed( in[140] ) ) - ( $signed( in[154] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_23;
always @( posedge clock ) begin
tree_23 <= ( $signed( in[17] ) ) - ( $signed( in[131] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_24;
always @( posedge clock ) begin
tree_24 <= ( $signed( in[62] ) ) + ( $signed( in[76] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_25;
always @( posedge clock ) begin
tree_25 <= ( $signed( in[15] ) ) + ( $signed( in[77] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_26;
always @( posedge clock ) begin
tree_26 <= ( $signed( in[132] ) ) + ( $signed( in[178] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_27;
always @( posedge clock ) begin
tree_27 <= ( $signed( in[122] ) ) + ( $signed( in[168] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_28;
always @( posedge clock ) begin
tree_28 <= ( $signed( in[151] ) ) + ( $signed( in[187] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_29;
always @( posedge clock ) begin
tree_29 <= ( $signed( in[114] ) ) + ( $signed( in[142] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_30;
always @( posedge clock ) begin
tree_30 <= ( $signed( in[24] ) ) - ( $signed( in[40] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_31;
always @( posedge clock ) begin
tree_31 <= ( $signed( in[47] ) ) - ( $signed( in[56] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_32;
always @( posedge clock ) begin
tree_32 <= ( $signed( in[74] ) ) + ( $signed( in[159] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_33;
always @( posedge clock ) begin
tree_33 <= ( $signed( in[148] ) ) + ( $signed( in[160] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_34;
always @( posedge clock ) begin
tree_34 <= ( $signed( in[38] ) ) + ( $signed( in[52] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_35;
always @( posedge clock ) begin
tree_35 <= ( $signed( in[126] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_36;
always @( posedge clock ) begin
tree_36 <= ( $signed( tree_35 ) ) + ( $signed( tree_19 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_37;
always @( posedge clock ) begin
tree_37 <= ( $signed( in[128] ) ) + ( $signed( in[186] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_38;
always @( posedge clock ) begin
tree_38 <= ( $signed( in[80] ) ) + ( $signed( in[83] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_39;
always @( posedge clock ) begin
tree_39 <= ( $signed( in[19] ) ) + ( $signed( in[59] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_40;
always @( posedge clock ) begin
tree_40 <= ( $signed( in[135] ) ) + ( $signed( in[180] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_41;
always @( posedge clock ) begin
tree_41 <= ( $signed( in[48] ) ) - ( $signed( in[140] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_42;
always @( posedge clock ) begin
tree_42 <= ( $signed( in[166] ) ) + ( $signed( in[188] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_43;
always @( posedge clock ) begin
tree_43 <= ( $signed( in[30] ) ) - ( $signed( in[44] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_44;
always @( posedge clock ) begin
tree_44 <= ( $signed( in[141] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_45;
always @( posedge clock ) begin
tree_45 <= ( $signed( tree_44 ) ) + ( $signed( tree_0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_46;
always @( posedge clock ) begin
tree_46 <= ( $signed( in[171] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_47;
always @( posedge clock ) begin
tree_47 <= ( $signed( tree_46 ) ) - ( $signed( tree_16 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_48;
always @( posedge clock ) begin
tree_48 <= ( $signed( in[85] ) ) - ( $signed( in[103] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_49;
always @( posedge clock ) begin
tree_49 <= ( $signed( in[142] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_50;
always @( posedge clock ) begin
tree_50 <= ( $signed( tree_49 ) ) - ( $signed( tree_2 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_51;
always @( posedge clock ) begin
tree_51 <= ( $signed( in[58] ) ) - ( $signed( in[174] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_52;
always @( posedge clock ) begin
tree_52 <= ( $signed( in[88] ) ) - ( $signed( in[173] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_53;
always @( posedge clock ) begin
tree_53 <= ( $signed( in[37] ) ) - ( $signed( in[109] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_54;
always @( posedge clock ) begin
tree_54 <= ( $signed( in[71] ) ) - ( $signed( in[106] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_55;
always @( posedge clock ) begin
tree_55 <= ( $signed( in[14] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_56;
always @( posedge clock ) begin
tree_56 <= ( $signed( tree_55 ) ) - ( $signed( tree_9 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_57;
always @( posedge clock ) begin
tree_57 <= ( $signed( in[81] ) ) + ( $signed( in[100] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_58;
always @( posedge clock ) begin
tree_58 <= ( $signed( in[84] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_59;
always @( posedge clock ) begin
tree_59 <= ( $signed( tree_58 ) ) + ( $signed( tree_18 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_60;
always @( posedge clock ) begin
tree_60 <= ( $signed( in[38] ) ) + ( $signed( in[79] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_61;
always @( posedge clock ) begin
tree_61 <= ( $signed( in[20] ) ) - ( $signed( in[33] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_62;
always @( posedge clock ) begin
tree_62 <= ( $signed( in[119] ) ) - ( $signed( in[173] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_63;
always @( posedge clock ) begin
tree_63 <= ( $signed( in[10] ) ) - ( $signed( in[61] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_64;
always @( posedge clock ) begin
tree_64 <= ( $signed( in[27] ) ) + ( $signed( in[56] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_65;
always @( posedge clock ) begin
tree_65 <= ( $signed( in[28] ) ) - ( $signed( in[91] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_66;
always @( posedge clock ) begin
tree_66 <= ( $signed( in[4] ) ) - ( $signed( in[77] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_67;
always @( posedge clock ) begin
tree_67 <= ( $signed( in[85] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_68;
always @( posedge clock ) begin
tree_68 <= ( $signed( tree_67 ) ) - ( $signed( tree_7 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_69;
always @( posedge clock ) begin
tree_69 <= ( $signed( in[116] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_70;
always @( posedge clock ) begin
tree_70 <= ( $signed( tree_69 ) ) - ( $signed( tree_6 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_71;
always @( posedge clock ) begin
tree_71 <= ( $signed( in[84] ) ) + ( $signed( in[167] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_72;
always @( posedge clock ) begin
tree_72 <= ( $signed( in[53] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_73;
always @( posedge clock ) begin
tree_73 <= ( $signed( tree_72 ) ) - ( $signed( tree_15 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_74;
always @( posedge clock ) begin
tree_74 <= ( $signed( in[25] ) ) + ( $signed( in[41] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_75;
always @( posedge clock ) begin
tree_75 <= ( $signed( in[89] ) ) + ( $signed( in[105] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_76;
always @( posedge clock ) begin
tree_76 <= ( $signed( in[127] ) ) + ( $signed( in[139] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_77;
always @( posedge clock ) begin
tree_77 <= ( $signed( in[60] ) ) - ( $signed( in[118] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_78;
always @( posedge clock ) begin
tree_78 <= ( $signed( in[132] ) ) - ( $signed( in[162] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_79;
always @( posedge clock ) begin
tree_79 <= ( $signed( in[93] ) ) + ( $signed( in[113] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_80;
always @( posedge clock ) begin
tree_80 <= ( $signed( in[72] ) ) + ( $signed( in[154] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_81;
always @( posedge clock ) begin
tree_81 <= ( $signed( in[16] ) ) - ( $signed( in[66] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_82;
always @( posedge clock ) begin
tree_82 <= ( $signed( in[65] ) ) - ( $signed( in[145] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_83;
always @( posedge clock ) begin
tree_83 <= ( $signed( in[146] ) ) - ( $signed( in[186] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_84;
always @( posedge clock ) begin
tree_84 <= ( $signed( in[86] ) ) + ( $signed( in[96] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_85;
always @( posedge clock ) begin
tree_85 <= ( $signed( in[100] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_86;
always @( posedge clock ) begin
tree_86 <= ( $signed( tree_85 ) ) + ( $signed( tree_32 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_87;
always @( posedge clock ) begin
tree_87 <= ( $signed( in[15] ) ) + ( $signed( in[63] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_88;
always @( posedge clock ) begin
tree_88 <= ( $signed( in[79] ) ) + ( $signed( in[97] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_89;
always @( posedge clock ) begin
tree_89 <= ( $signed( in[155] ) ) + ( $signed( in[179] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_90;
always @( posedge clock ) begin
tree_90 <= ( $signed( in[93] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_91;
always @( posedge clock ) begin
tree_91 <= ( $signed( tree_90 ) ) - ( $signed( tree_16 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_92;
always @( posedge clock ) begin
tree_92 <= ( $signed( in[135] ) ) - ( $signed( in[169] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_93;
always @( posedge clock ) begin
tree_93 <= ( $signed( in[6] ) ) + ( $signed( in[177] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_94;
always @( posedge clock ) begin
tree_94 <= ( $signed( in[82] ) ) - ( $signed( in[145] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_95;
always @( posedge clock ) begin
tree_95 <= ( $signed( in[136] ) ) - ( $signed( in[185] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_96;
always @( posedge clock ) begin
tree_96 <= ( $signed( in[131] ) ) + ( $signed( in[149] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_97;
always @( posedge clock ) begin
tree_97 <= ( $signed( in[55] ) ) - ( $signed( in[116] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_98;
always @( posedge clock ) begin
tree_98 <= ( $signed( tree_28 ) ) - ( $signed( tree_18 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_99;
always @( posedge clock ) begin
tree_99 <= ( $signed( in[30] ) ) + ( $signed( in[50] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_100;
always @( posedge clock ) begin
tree_100 <= ( $signed( in[14] ) ) + ( $signed( in[20] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_101;
always @( posedge clock ) begin
tree_101 <= ( $signed( in[2] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_102;
always @( posedge clock ) begin
tree_102 <= ( $signed( tree_101 ) ) - ( $signed( tree_21 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_103;
always @( posedge clock ) begin
tree_103 <= ( $signed( in[24] ) ) + ( $signed( in[164] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_104;
always @( posedge clock ) begin
tree_104 <= ( $signed( in[142] ) ) + ( $signed( in[172] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_105;
always @( posedge clock ) begin
tree_105 <= ( $signed( in[184] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_106;
always @( posedge clock ) begin
tree_106 <= ( $signed( tree_105 ) ) + ( $signed( tree_20 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_107;
always @( posedge clock ) begin
tree_107 <= ( $signed( in[62] ) ) - ( $signed( in[66] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_108;
always @( posedge clock ) begin
tree_108 <= ( $signed( in[5] ) ) - ( $signed( in[70] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_109;
always @( posedge clock ) begin
tree_109 <= ( $signed( in[35] ) ) - ( $signed( in[87] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_110;
always @( posedge clock ) begin
tree_110 <= ( $signed( in[121] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_111;
always @( posedge clock ) begin
tree_111 <= ( $signed( tree_110 ) ) - ( $signed( tree_64 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_112;
always @( posedge clock ) begin
tree_112 <= ( $signed( in[7] ) ) - ( $signed( in[86] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_113;
always @( posedge clock ) begin
tree_113 <= ( $signed( in[134] ) ) + ( $signed( in[176] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_114;
always @( posedge clock ) begin
tree_114 <= ( $signed( in[90] ) ) - ( $signed( in[120] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_115;
always @( posedge clock ) begin
tree_115 <= ( $signed( in[110] ) ) + ( $signed( in[150] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_116;
always @( posedge clock ) begin
tree_116 <= ( $signed( in[167] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_117;
always @( posedge clock ) begin
tree_117 <= ( $signed( tree_116 ) ) + ( $signed( tree_0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_118;
always @( posedge clock ) begin
tree_118 <= ( $signed( in[131] ) ) - ( $signed( in[172] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_119;
always @( posedge clock ) begin
tree_119 <= ( $signed( in[10] ) ) - ( $signed( in[52] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_120;
always @( posedge clock ) begin
tree_120 <= ( $signed( in[49] ) ) - ( $signed( in[170] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_121;
always @( posedge clock ) begin
tree_121 <= ( $signed( in[45] ) ) - ( $signed( in[88] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_122;
always @( posedge clock ) begin
tree_122 <= ( $signed( in[116] ) ) - ( $signed( in[129] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_123;
always @( posedge clock ) begin
tree_123 <= ( $signed( in[97] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_124;
always @( posedge clock ) begin
tree_124 <= ( $signed( tree_123 ) ) - ( $signed( tree_40 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_125;
always @( posedge clock ) begin
tree_125 <= ( $signed( in[30] ) ) - ( $signed( in[46] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_126;
always @( posedge clock ) begin
tree_126 <= ( $signed( in[84] ) ) - ( $signed( in[183] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_127;
always @( posedge clock ) begin
tree_127 <= ( $signed( in[152] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_128;
always @( posedge clock ) begin
tree_128 <= ( $signed( tree_127 ) ) - ( $signed( tree_11 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_129;
always @( posedge clock ) begin
tree_129 <= ( $signed( in[11] ) ) + ( $signed( in[78] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_130;
always @( posedge clock ) begin
tree_130 <= ( $signed( in[73] ) ) + ( $signed( in[158] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_131;
always @( posedge clock ) begin
tree_131 <= ( $signed( in[126] ) ) + ( $signed( in[173] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_132;
always @( posedge clock ) begin
tree_132 <= ( $signed( in[9] ) ) - ( $signed( in[159] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_133;
always @( posedge clock ) begin
tree_133 <= ( $signed( in[67] ) ) - ( $signed( in[113] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_134;
always @( posedge clock ) begin
tree_134 <= ( $signed( in[57] ) ) - ( $signed( in[82] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_135;
always @( posedge clock ) begin
tree_135 <= ( $signed( in[36] ) ) + ( $signed( in[49] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_136;
always @( posedge clock ) begin
tree_136 <= ( $signed( in[157] ) ) + ( $signed( in[168] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_137;
always @( posedge clock ) begin
tree_137 <= ( $signed( in[48] ) ) - ( $signed( in[166] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_138;
always @( posedge clock ) begin
tree_138 <= ( $signed( in[43] ) ) - ( $signed( in[69] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_139;
always @( posedge clock ) begin
tree_139 <= ( $signed( in[13] ) ) + ( $signed( in[44] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_140;
always @( posedge clock ) begin
tree_140 <= ( $signed( in[99] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_141;
always @( posedge clock ) begin
tree_141 <= ( $signed( tree_140 ) ) - ( $signed( tree_22 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_142;
always @( posedge clock ) begin
tree_142 <= ( $signed( in[55] ) ) - ( $signed( in[63] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_143;
always @( posedge clock ) begin
tree_143 <= ( $signed( in[17] ) ) - ( $signed( in[60] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_144;
always @( posedge clock ) begin
tree_144 <= ( $signed( tree_21 ) ) - ( $signed( tree_122 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_145;
always @( posedge clock ) begin
tree_145 <= ( $signed( in[5] ) ) - ( $signed( in[99] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_146;
always @( posedge clock ) begin
tree_146 <= ( $signed( in[75] ) ) - ( $signed( in[176] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_147;
always @( posedge clock ) begin
tree_147 <= ( $signed( in[3] ) ) + ( $signed( in[11] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_148;
always @( posedge clock ) begin
tree_148 <= ( $signed( in[66] ) ) - ( $signed( in[77] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_149;
always @( posedge clock ) begin
tree_149 <= ( $signed( in[37] ) ) - ( $signed( in[126] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_150;
always @( posedge clock ) begin
tree_150 <= ( $signed( in[114] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_151;
always @( posedge clock ) begin
tree_151 <= ( $signed( tree_150 ) ) - ( $signed( tree_74 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_152;
always @( posedge clock ) begin
tree_152 <= ( $signed( in[12] ) ) + ( $signed( in[134] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_153;
always @( posedge clock ) begin
tree_153 <= ( $signed( in[112] ) ) + ( $signed( in[125] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_154;
always @( posedge clock ) begin
tree_154 <= ( $signed( in[85] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_155;
always @( posedge clock ) begin
tree_155 <= ( $signed( tree_154 ) ) - ( $signed( tree_3 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_156;
always @( posedge clock ) begin
tree_156 <= ( $signed( in[191] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_157;
always @( posedge clock ) begin
tree_157 <= ( $signed( tree_156 ) ) - ( $signed( tree_41 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_158;
always @( posedge clock ) begin
tree_158 <= ( $signed( in[183] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_159;
always @( posedge clock ) begin
tree_159 <= ( $signed( tree_158 ) ) + ( $signed( tree_26 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_160;
always @( posedge clock ) begin
tree_160 <= ( $signed( tree_32 ) ) - ( $signed( tree_92 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_161;
always @( posedge clock ) begin
tree_161 <= ( $signed( in[65] ) ) - ( $signed( in[103] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_162;
always @( posedge clock ) begin
tree_162 <= ( $signed( in[29] ) ) + ( $signed( in[138] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_163;
always @( posedge clock ) begin
tree_163 <= ( $signed( in[108] ) ) - ( $signed( in[139] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_164;
always @( posedge clock ) begin
tree_164 <= ( $signed( in[0] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_165;
always @( posedge clock ) begin
tree_165 <= ( $signed( tree_164 ) ) + ( $signed( tree_139 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_166;
always @( posedge clock ) begin
tree_166 <= ( $signed( in[1] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_167;
always @( posedge clock ) begin
tree_167 <= ( $signed( tree_166 ) ) + ( $signed( tree_30 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_168;
always @( posedge clock ) begin
tree_168 <= ( $signed( in[32] ) ) - ( $signed( in[157] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_169;
always @( posedge clock ) begin
tree_169 <= ( $signed( in[43] ) ) - ( $signed( in[154] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_170;
always @( posedge clock ) begin
tree_170 <= ( $signed( in[46] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_171;
always @( posedge clock ) begin
tree_171 <= ( $signed( tree_170 ) ) - ( $signed( tree_81 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_172;
always @( posedge clock ) begin
tree_172 <= ( $signed( in[104] ) ) + ( $signed( in[165] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_173;
always @( posedge clock ) begin
tree_173 <= ( $signed( in[164] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_174;
always @( posedge clock ) begin
tree_174 <= ( $signed( tree_173 ) ) - ( $signed( tree_79 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_175;
always @( posedge clock ) begin
tree_175 <= ( $signed( in[172] ) ) - ( $signed( in[178] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_176;
always @( posedge clock ) begin
tree_176 <= ( $signed( in[74] ) ) + ( $signed( in[110] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_177;
always @( posedge clock ) begin
tree_177 <= ( $signed( in[24] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_178;
always @( posedge clock ) begin
tree_178 <= ( $signed( tree_177 ) ) + ( $signed( tree_78 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_179;
always @( posedge clock ) begin
tree_179 <= ( $signed( in[51] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_180;
always @( posedge clock ) begin
tree_180 <= ( $signed( tree_179 ) ) + ( $signed( tree_42 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_181;
always @( posedge clock ) begin
tree_181 <= ( $signed( in[38] ) ) - ( $signed( in[103] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_182;
always @( posedge clock ) begin
tree_182 <= ( $signed( in[190] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_183;
always @( posedge clock ) begin
tree_183 <= ( $signed( tree_182 ) ) - ( $signed( tree_65 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_184;
always @( posedge clock ) begin
tree_184 <= ( $signed( in[182] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_185;
always @( posedge clock ) begin
tree_185 <= ( $signed( tree_184 ) ) - ( $signed( tree_9 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_186;
always @( posedge clock ) begin
tree_186 <= ( $signed( in[73] ) ) - ( $signed( in[134] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_187;
always @( posedge clock ) begin
tree_187 <= ( $signed( in[98] ) ) + ( $signed( in[103] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_188;
always @( posedge clock ) begin
tree_188 <= ( $signed( in[5] ) ) - ( $signed( in[188] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_189;
always @( posedge clock ) begin
tree_189 <= ( $signed( in[1] ) ) - ( $signed( in[45] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_190;
always @( posedge clock ) begin
tree_190 <= ( $signed( in[76] ) ) - ( $signed( in[127] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_191;
always @( posedge clock ) begin
tree_191 <= ( $signed( in[95] ) ) - ( $signed( in[136] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_192;
always @( posedge clock ) begin
tree_192 <= ( $signed( in[6] ) ) - ( $signed( in[89] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_193;
always @( posedge clock ) begin
tree_193 <= ( $signed( in[27] ) ) - ( $signed( in[137] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_194;
always @( posedge clock ) begin
tree_194 <= ( $signed( in[49] ) ) - ( $signed( in[63] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_195;
always @( posedge clock ) begin
tree_195 <= ( $signed( in[14] ) ) + ( $signed( in[65] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_196;
always @( posedge clock ) begin
tree_196 <= ( $signed( in[10] ) ) - ( $signed( in[99] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_197;
always @( posedge clock ) begin
tree_197 <= ( $signed( in[147] ) ) + ( $signed( in[157] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_198;
always @( posedge clock ) begin
tree_198 <= ( $signed( in[32] ) ) - ( $signed( in[156] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_199;
always @( posedge clock ) begin
tree_199 <= ( $signed( in[82] ) ) + ( $signed( in[85] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_200;
always @( posedge clock ) begin
tree_200 <= ( $signed( in[70] ) ) + ( $signed( in[79] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_201;
always @( posedge clock ) begin
tree_201 <= ( $signed( in[116] ) ) + ( $signed( in[153] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_202;
always @( posedge clock ) begin
tree_202 <= ( $signed( in[7] ) ) - ( $signed( in[33] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_203;
always @( posedge clock ) begin
tree_203 <= ( $signed( in[81] ) ) - ( $signed( in[85] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_204;
always @( posedge clock ) begin
tree_204 <= ( $signed( in[3] ) ) - ( $signed( in[36] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_205;
always @( posedge clock ) begin
tree_205 <= ( $signed( in[115] ) ) + ( $signed( in[139] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_206;
always @( posedge clock ) begin
tree_206 <= ( $signed( in[18] ) ) - ( $signed( in[142] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_207;
always @( posedge clock ) begin
tree_207 <= ( $signed( in[114] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_208;
always @( posedge clock ) begin
tree_208 <= ( $signed( tree_207 ) ) - ( $signed( tree_10 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_209;
always @( posedge clock ) begin
tree_209 <= ( $signed( in[22] ) ) - ( $signed( in[29] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_210;
always @( posedge clock ) begin
tree_210 <= ( $signed( in[23] ) ) + ( $signed( in[59] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_211;
always @( posedge clock ) begin
tree_211 <= ( $signed( in[143] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_212;
always @( posedge clock ) begin
tree_212 <= ( $signed( tree_211 ) ) + ( $signed( tree_7 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_213;
always @( posedge clock ) begin
tree_213 <= ( $signed( in[2] ) ) + ( $signed( in[46] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_214;
always @( posedge clock ) begin
tree_214 <= ( $signed( in[68] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_215;
always @( posedge clock ) begin
tree_215 <= ( $signed( tree_214 ) ) - ( $signed( tree_89 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_216;
always @( posedge clock ) begin
tree_216 <= ( $signed( in[20] ) ) + ( $signed( in[31] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_217;
always @( posedge clock ) begin
tree_217 <= ( $signed( in[4] ) ) - ( $signed( in[56] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_218;
always @( posedge clock ) begin
tree_218 <= ( $signed( tree_142 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_219;
always @( posedge clock ) begin
tree_219 <=  - ( $signed( tree_218 ) ) + ( $signed( tree_36 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_220;
always @( posedge clock ) begin
tree_220 <= ( $signed( in[98] ) ) - ( $signed( in[183] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_221;
always @( posedge clock ) begin
tree_221 <= ( $signed( in[53] ) ) - ( $signed( in[96] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_222;
always @( posedge clock ) begin
tree_222 <= ( $signed( in[45] ) ) + ( $signed( in[174] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_223;
always @( posedge clock ) begin
tree_223 <= ( $signed( in[51] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_224;
always @( posedge clock ) begin
tree_224 <= ( $signed( tree_223 ) ) - ( $signed( tree_88 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_225;
always @( posedge clock ) begin
tree_225 <= ( $signed( in[8] ) ) + ( $signed( in[44] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_226;
always @( posedge clock ) begin
tree_226 <= ( $signed( in[3] ) ) - ( $signed( in[55] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_227;
always @( posedge clock ) begin
tree_227 <= ( $signed( in[155] ) ) - ( $signed( in[168] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_228;
always @( posedge clock ) begin
tree_228 <= ( $signed( in[84] ) ) - ( $signed( in[128] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_229;
always @( posedge clock ) begin
tree_229 <= ( $signed( in[12] ) ) - ( $signed( in[18] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_230;
always @( posedge clock ) begin
tree_230 <= ( $signed( in[101] ) ) - ( $signed( in[149] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_231;
always @( posedge clock ) begin
tree_231 <= ( $signed( in[33] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_232;
always @( posedge clock ) begin
tree_232 <= ( $signed( tree_231 ) ) - ( $signed( tree_74 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_233;
always @( posedge clock ) begin
tree_233 <= ( $signed( in[47] ) ) - ( $signed( in[94] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_234;
always @( posedge clock ) begin
tree_234 <= ( $signed( in[108] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_235;
always @( posedge clock ) begin
tree_235 <= ( $signed( tree_234 ) ) - ( $signed( tree_16 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_236;
always @( posedge clock ) begin
tree_236 <= ( $signed( in[112] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_237;
always @( posedge clock ) begin
tree_237 <= ( $signed( tree_236 ) ) - ( $signed( tree_161 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_238;
always @( posedge clock ) begin
tree_238 <= ( $signed( in[98] ) ) + ( $signed( in[130] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_239;
always @( posedge clock ) begin
tree_239 <= ( $signed( tree_88 ) ) + ( $signed( tree_119 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_240;
always @( posedge clock ) begin
tree_240 <= ( $signed( tree_13 ) ) - ( $signed( tree_186 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_241;
always @( posedge clock ) begin
tree_241 <= ( $signed( in[82] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_242;
always @( posedge clock ) begin
tree_242 <= ( $signed( tree_241 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_243;
always @( posedge clock ) begin
tree_243 <= ( $signed( tree_242 ) ) + ( $signed( tree_86 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_244;
always @( posedge clock ) begin
tree_244 <= ( $signed( in[143] ) ) - ( $signed( in[151] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_245;
always @( posedge clock ) begin
tree_245 <= ( $signed( in[24] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_246;
always @( posedge clock ) begin
tree_246 <= ( $signed( tree_245 ) ) - ( $signed( tree_7 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_247;
always @( posedge clock ) begin
tree_247 <= ( $signed( in[111] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_248;
always @( posedge clock ) begin
tree_248 <= ( $signed( tree_247 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_249;
always @( posedge clock ) begin
tree_249 <= ( $signed( tree_248 ) ) + ( $signed( tree_159 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_250;
always @( posedge clock ) begin
tree_250 <= ( $signed( in[15] ) ) - ( $signed( in[159] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_251;
always @( posedge clock ) begin
tree_251 <= ( $signed( in[62] ) ) - ( $signed( in[138] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_252;
always @( posedge clock ) begin
tree_252 <= ( $signed( in[186] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_253;
always @( posedge clock ) begin
tree_253 <= ( $signed( tree_252 ) ) - ( $signed( tree_82 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_254;
always @( posedge clock ) begin
tree_254 <= ( $signed( in[20] ) ) - ( $signed( in[161] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_255;
always @( posedge clock ) begin
tree_255 <= ( $signed( in[67] ) ) - ( $signed( in[78] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_256;
always @( posedge clock ) begin
tree_256 <= ( $signed( in[125] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_257;
always @( posedge clock ) begin
tree_257 <= ( $signed( tree_256 ) ) - ( $signed( tree_74 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_258;
always @( posedge clock ) begin
tree_258 <= ( $signed( in[4] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_259;
always @( posedge clock ) begin
tree_259 <= ( $signed( tree_258 ) ) + ( $signed( tree_21 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_260;
always @( posedge clock ) begin
tree_260 <= ( $signed( in[17] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_261;
always @( posedge clock ) begin
tree_261 <= ( $signed( tree_260 ) ) - ( $signed( tree_96 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_262;
always @( posedge clock ) begin
tree_262 <= ( $signed( in[16] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_263;
always @( posedge clock ) begin
tree_263 <= ( $signed( tree_262 ) ) - ( $signed( tree_63 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_264;
always @( posedge clock ) begin
tree_264 <= ( $signed( in[51] ) ) - ( $signed( in[170] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_265;
always @( posedge clock ) begin
tree_265 <= ( $signed( in[19] ) ) - ( $signed( in[75] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_266;
always @( posedge clock ) begin
tree_266 <= ( $signed( in[16] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_267;
always @( posedge clock ) begin
tree_267 <= ( $signed( tree_266 ) ) - ( $signed( tree_4 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_268;
always @( posedge clock ) begin
tree_268 <= ( $signed( in[44] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_269;
always @( posedge clock ) begin
tree_269 <= ( $signed( tree_268 ) ) - ( $signed( tree_34 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_270;
always @( posedge clock ) begin
tree_270 <= ( $signed( in[33] ) ) - ( $signed( in[146] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_271;
always @( posedge clock ) begin
tree_271 <= ( $signed( in[13] ) ) - ( $signed( in[139] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_272;
always @( posedge clock ) begin
tree_272 <= ( $signed( in[35] ) ) - ( $signed( in[124] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_273;
always @( posedge clock ) begin
tree_273 <= ( $signed( in[58] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_274;
always @( posedge clock ) begin
tree_274 <= ( $signed( tree_273 ) ) + ( $signed( tree_210 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_275;
always @( posedge clock ) begin
tree_275 <= ( $signed( in[57] ) ) - ( $signed( in[86] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_276;
always @( posedge clock ) begin
tree_276 <= ( $signed( in[6] ) ) + ( $signed( in[68] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_277;
always @( posedge clock ) begin
tree_277 <= ( $signed( in[98] ) ) + ( $signed( in[175] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_278;
always @( posedge clock ) begin
tree_278 <= ( $signed( in[40] ) ) - ( $signed( in[62] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_279;
always @( posedge clock ) begin
tree_279 <= ( $signed( tree_57 ) ) - ( $signed( tree_189 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_280;
always @( posedge clock ) begin
tree_280 <= ( $signed( in[61] ) ) + ( $signed( in[189] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_281;
always @( posedge clock ) begin
tree_281 <= ( $signed( in[68] ) ) + ( $signed( in[153] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_282;
always @( posedge clock ) begin
tree_282 <= ( $signed( tree_147 ) ) + ( $signed( tree_188 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_283;
always @( posedge clock ) begin
tree_283 <= ( $signed( tree_146 ) ) - ( $signed( tree_22 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_284;
always @( posedge clock ) begin
tree_284 <= ( $signed( in[102] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_285;
always @( posedge clock ) begin
tree_285 <= ( $signed( tree_284 ) ) - ( $signed( tree_210 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_286;
always @( posedge clock ) begin
tree_286 <= ( $signed( in[166] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_287;
always @( posedge clock ) begin
tree_287 <= ( $signed( tree_286 ) ) - ( $signed( tree_27 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_288;
always @( posedge clock ) begin
tree_288 <= ( $signed( in[3] ) ) + ( $signed( in[149] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_289;
always @( posedge clock ) begin
tree_289 <= ( $signed( in[41] ) ) - ( $signed( in[140] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_290;
always @( posedge clock ) begin
tree_290 <= ( $signed( in[23] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_291;
always @( posedge clock ) begin
tree_291 <= ( $signed( tree_290 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_292;
always @( posedge clock ) begin
tree_292 <= ( $signed( tree_291 ) ) - ( $signed( tree_215 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_293;
always @( posedge clock ) begin
tree_293 <= ( $signed( in[118] ) ) + ( $signed( in[145] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_294;
always @( posedge clock ) begin
tree_294 <= ( $signed( in[8] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_295;
always @( posedge clock ) begin
tree_295 <= ( $signed( tree_294 ) ) - ( $signed( tree_53 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_296;
always @( posedge clock ) begin
tree_296 <= ( $signed( in[93] ) ) - ( $signed( in[151] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_297;
always @( posedge clock ) begin
tree_297 <= ( $signed( in[165] ) ) - ( $signed( in[175] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_298;
always @( posedge clock ) begin
tree_298 <= ( $signed( in[28] ) ) - ( $signed( in[158] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_299;
always @( posedge clock ) begin
tree_299 <= ( $signed( tree_135 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_300;
always @( posedge clock ) begin
tree_300 <= ( $signed( tree_299 ) ) - ( $signed( tree_117 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_301;
always @( posedge clock ) begin
tree_301 <= ( $signed( in[84] ) ) + ( $signed( in[182] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_302;
always @( posedge clock ) begin
tree_302 <= ( $signed( in[98] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_303;
always @( posedge clock ) begin
tree_303 <= ( $signed( tree_302 ) ) + ( $signed( tree_76 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_304;
always @( posedge clock ) begin
tree_304 <= ( $signed( in[26] ) ) - ( $signed( in[177] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_305;
always @( posedge clock ) begin
tree_305 <= ( $signed( in[188] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_306;
always @( posedge clock ) begin
tree_306 <= ( $signed( tree_305 ) ) - ( $signed( tree_195 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_307;
always @( posedge clock ) begin
tree_307 <= ( $signed( in[109] ) ) + ( $signed( in[162] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_308;
always @( posedge clock ) begin
tree_308 <= ( $signed( in[14] ) ) - ( $signed( in[93] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_309;
always @( posedge clock ) begin
tree_309 <= ( $signed( in[149] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_310;
always @( posedge clock ) begin
tree_310 <= ( $signed( tree_309 ) ) - ( $signed( tree_27 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_311;
always @( posedge clock ) begin
tree_311 <= ( $signed( tree_14 ) ) - ( $signed( tree_80 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_312;
always @( posedge clock ) begin
tree_312 <= ( $signed( in[12] ) ) + ( $signed( in[140] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_313;
always @( posedge clock ) begin
tree_313 <= ( $signed( in[19] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_314;
always @( posedge clock ) begin
tree_314 <= ( $signed( tree_313 ) ) - ( $signed( tree_71 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_315;
always @( posedge clock ) begin
tree_315 <= ( $signed( in[123] ) ) - ( $signed( in[185] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_316;
always @( posedge clock ) begin
tree_316 <= ( $signed( in[136] ) ) + ( $signed( in[146] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_317;
always @( posedge clock ) begin
tree_317 <= ( $signed( in[147] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_318;
always @( posedge clock ) begin
tree_318 <= ( $signed( tree_317 ) ) - ( $signed( tree_103 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_319;
always @( posedge clock ) begin
tree_319 <= ( $signed( in[90] ) ) - ( $signed( in[190] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_320;
always @( posedge clock ) begin
tree_320 <= ( $signed( in[104] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_321;
always @( posedge clock ) begin
tree_321 <= ( $signed( tree_320 ) ) - ( $signed( tree_87 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_322;
always @( posedge clock ) begin
tree_322 <= ( $signed( in[102] ) ) + ( $signed( in[191] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_323;
always @( posedge clock ) begin
tree_323 <= ( $signed( in[52] ) ) - ( $signed( in[152] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_324;
always @( posedge clock ) begin
tree_324 <= ( $signed( in[60] ) ) - ( $signed( in[106] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_325;
always @( posedge clock ) begin
tree_325 <= ( $signed( in[91] ) ) + ( $signed( in[171] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_326;
always @( posedge clock ) begin
tree_326 <= ( $signed( in[24] ) ) - ( $signed( in[143] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_327;
always @( posedge clock ) begin
tree_327 <= ( $signed( in[111] ) ) - ( $signed( in[153] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_328;
always @( posedge clock ) begin
tree_328 <= ( $signed( in[25] ) ) - ( $signed( in[120] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_329;
always @( posedge clock ) begin
tree_329 <= ( $signed( in[96] ) ) + ( $signed( in[189] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_330;
always @( posedge clock ) begin
tree_330 <= ( $signed( in[13] ) ) - ( $signed( in[129] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_331;
always @( posedge clock ) begin
tree_331 <= ( $signed( in[14] ) ) - ( $signed( in[16] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_332;
always @( posedge clock ) begin
tree_332 <= ( $signed( in[53] ) ) - ( $signed( in[69] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_333;
always @( posedge clock ) begin
tree_333 <= ( $signed( in[19] ) ) + ( $signed( in[77] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_334;
always @( posedge clock ) begin
tree_334 <= ( $signed( in[107] ) ) + ( $signed( in[137] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_335;
always @( posedge clock ) begin
tree_335 <= ( $signed( in[71] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_336;
always @( posedge clock ) begin
tree_336 <= ( $signed( tree_335 ) ) - ( $signed( tree_202 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_337;
always @( posedge clock ) begin
tree_337 <= ( $signed( in[94] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_338;
always @( posedge clock ) begin
tree_338 <= ( $signed( tree_337 ) ) - ( $signed( tree_17 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_339;
always @( posedge clock ) begin
tree_339 <= ( $signed( in[47] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_340;
always @( posedge clock ) begin
tree_340 <= ( $signed( tree_339 ) ) + ( $signed( tree_187 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_341;
always @( posedge clock ) begin
tree_341 <= ( $signed( in[1] ) ) - ( $signed( in[107] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_342;
always @( posedge clock ) begin
tree_342 <= ( $signed( in[6] ) ) - ( $signed( in[22] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_343;
always @( posedge clock ) begin
tree_343 <= ( $signed( in[50] ) ) - ( $signed( in[118] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_344;
always @( posedge clock ) begin
tree_344 <= ( $signed( in[78] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_345;
always @( posedge clock ) begin
tree_345 <= ( $signed( tree_344 ) ) - ( $signed( tree_28 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_346;
always @( posedge clock ) begin
tree_346 <= ( $signed( in[37] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_347;
always @( posedge clock ) begin
tree_347 <= ( $signed( tree_346 ) ) - ( $signed( tree_29 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_348;
always @( posedge clock ) begin
tree_348 <= ( $signed( in[61] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_349;
always @( posedge clock ) begin
tree_349 <= ( $signed( tree_348 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_350;
always @( posedge clock ) begin
tree_350 <= ( $signed( tree_349 ) ) - ( $signed( tree_106 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_351;
always @( posedge clock ) begin
tree_351 <= ( $signed( in[109] ) ) - ( $signed( in[134] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_352;
always @( posedge clock ) begin
tree_352 <= ( $signed( in[34] ) ) - ( $signed( in[165] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_353;
always @( posedge clock ) begin
tree_353 <= ( $signed( in[105] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_354;
always @( posedge clock ) begin
tree_354 <= ( $signed( tree_353 ) ) + ( $signed( tree_187 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_355;
always @( posedge clock ) begin
tree_355 <= ( $signed( in[86] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_356;
always @( posedge clock ) begin
tree_356 <= ( $signed( tree_355 ) ) - ( $signed( tree_143 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_357;
always @( posedge clock ) begin
tree_357 <= ( $signed( in[117] ) ) - ( $signed( in[122] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_358;
always @( posedge clock ) begin
tree_358 <= ( $signed( in[9] ) ) - ( $signed( in[64] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_359;
always @( posedge clock ) begin
tree_359 <= ( $signed( tree_146 ) ) - ( $signed( tree_40 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_360;
always @( posedge clock ) begin
tree_360 <= ( $signed( in[74] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_361;
always @( posedge clock ) begin
tree_361 <= ( $signed( tree_360 ) ) - ( $signed( tree_38 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_362;
always @( posedge clock ) begin
tree_362 <= ( $signed( in[34] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_363;
always @( posedge clock ) begin
tree_363 <= ( $signed( tree_362 ) ) - ( $signed( tree_188 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_364;
always @( posedge clock ) begin
tree_364 <= ( $signed( in[108] ) ) + ( $signed( in[173] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_365;
always @( posedge clock ) begin
tree_365 <= ( $signed( in[128] ) ) - ( $signed( in[175] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_366;
always @( posedge clock ) begin
tree_366 <= ( $signed( in[44] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_367;
always @( posedge clock ) begin
tree_367 <= ( $signed( tree_366 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_368;
always @( posedge clock ) begin
tree_368 <= ( $signed( tree_367 ) ) - ( $signed( tree_356 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_369;
always @( posedge clock ) begin
tree_369 <= ( $signed( in[65] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_370;
always @( posedge clock ) begin
tree_370 <= ( $signed( tree_369 ) ) - ( $signed( tree_312 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_371;
always @( posedge clock ) begin
tree_371 <= ( $signed( in[112] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_372;
always @( posedge clock ) begin
tree_372 <= ( $signed( tree_371 ) ) - ( $signed( tree_198 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_373;
always @( posedge clock ) begin
tree_373 <= ( $signed( tree_322 ) ) - ( $signed( tree_118 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_374;
always @( posedge clock ) begin
tree_374 <= ( $signed( in[150] ) ) - ( $signed( in[154] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_375;
always @( posedge clock ) begin
tree_375 <= ( $signed( tree_216 ) ) + ( $signed( tree_276 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_376;
always @( posedge clock ) begin
tree_376 <= ( $signed( in[27] ) ) - ( $signed( in[112] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_377;
always @( posedge clock ) begin
tree_377 <= ( $signed( tree_26 ) ) + ( $signed( tree_33 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_378;
always @( posedge clock ) begin
tree_378 <= ( $signed( in[38] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_379;
always @( posedge clock ) begin
tree_379 <= ( $signed( tree_378 ) ) - ( $signed( tree_152 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_380;
always @( posedge clock ) begin
tree_380 <= ( $signed( in[26] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_381;
always @( posedge clock ) begin
tree_381 <= ( $signed( tree_380 ) ) - ( $signed( tree_32 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_382;
always @( posedge clock ) begin
tree_382 <= ( $signed( in[113] ) ) + ( $signed( in[181] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_383;
always @( posedge clock ) begin
tree_383 <= ( $signed( in[126] ) ) - ( $signed( in[154] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_384;
always @( posedge clock ) begin
tree_384 <= ( $signed( tree_47 ) ) - ( $signed( tree_208 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_385;
always @( posedge clock ) begin
tree_385 <= ( $signed( in[101] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_386;
always @( posedge clock ) begin
tree_386 <= ( $signed( tree_385 ) ) + ( $signed( tree_280 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_387;
always @( posedge clock ) begin
tree_387 <= ( $signed( in[50] ) ) - ( $signed( in[151] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_388;
always @( posedge clock ) begin
tree_388 <= ( $signed( in[124] ) ) - ( $signed( in[133] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_389;
always @( posedge clock ) begin
tree_389 <= ( $signed( in[120] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_390;
always @( posedge clock ) begin
tree_390 <= ( $signed( tree_389 ) ) - ( $signed( tree_332 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_391;
always @( posedge clock ) begin
tree_391 <= ( $signed( in[21] ) ) - ( $signed( in[77] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_392;
always @( posedge clock ) begin
tree_392 <= ( $signed( in[127] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_393;
always @( posedge clock ) begin
tree_393 <= ( $signed( tree_392 ) ) - ( $signed( tree_162 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_394;
always @( posedge clock ) begin
tree_394 <= ( $signed( in[7] ) ) + ( $signed( in[45] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_395;
always @( posedge clock ) begin
tree_395 <= ( $signed( in[141] ) ) - ( $signed( in[174] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_396;
always @( posedge clock ) begin
tree_396 <= ( $signed( in[102] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_397;
always @( posedge clock ) begin
tree_397 <= ( $signed( tree_396 ) ) - ( $signed( tree_53 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_398;
always @( posedge clock ) begin
tree_398 <= ( $signed( in[36] ) ) - ( $signed( in[152] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_399;
always @( posedge clock ) begin
tree_399 <= ( $signed( tree_267 ) ) - ( $signed( tree_174 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_400;
always @( posedge clock ) begin
tree_400 <= ( $signed( in[135] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_401;
always @( posedge clock ) begin
tree_401 <= ( $signed( tree_400 ) ) - ( $signed( tree_6 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_402;
always @( posedge clock ) begin
tree_402 <= ( $signed( tree_78 ) ) + ( $signed( tree_130 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_403;
always @( posedge clock ) begin
tree_403 <= ( $signed( in[34] ) ) - ( $signed( in[48] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_404;
always @( posedge clock ) begin
tree_404 <= ( $signed( in[64] ) ) - ( $signed( in[144] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_405;
always @( posedge clock ) begin
tree_405 <= ( $signed( tree_63 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_406;
always @( posedge clock ) begin
tree_406 <= ( $signed( tree_405 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_407;
always @( posedge clock ) begin
tree_407 <= ( $signed( tree_406 ) ) - ( $signed( tree_292 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_408;
always @( posedge clock ) begin
tree_408 <= ( $signed( in[7] ) ) - ( $signed( in[184] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_409;
always @( posedge clock ) begin
tree_409 <= ( $signed( in[103] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_410;
always @( posedge clock ) begin
tree_410 <= ( $signed( tree_409 ) ) - ( $signed( tree_322 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_411;
always @( posedge clock ) begin
tree_411 <= ( $signed( in[83] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_412;
always @( posedge clock ) begin
tree_412 <= ( $signed( tree_411 ) ) + ( $signed( tree_143 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_413;
always @( posedge clock ) begin
tree_413 <= ( $signed( in[20] ) ) - ( $signed( in[158] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_414;
always @( posedge clock ) begin
tree_414 <= ( $signed( in[52] ) ) - ( $signed( in[167] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_415;
always @( posedge clock ) begin
tree_415 <= ( $signed( in[73] ) ) - ( $signed( in[181] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_416;
always @( posedge clock ) begin
tree_416 <= ( $signed( in[0] ) ) + ( $signed( in[171] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_417;
always @( posedge clock ) begin
tree_417 <= ( $signed( in[156] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_418;
always @( posedge clock ) begin
tree_418 <= ( $signed( tree_417 ) ) - ( $signed( tree_87 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_419;
always @( posedge clock ) begin
tree_419 <= ( $signed( in[8] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_420;
always @( posedge clock ) begin
tree_420 <= ( $signed( tree_419 ) ) - ( $signed( tree_78 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_421;
always @( posedge clock ) begin
tree_421 <= ( $signed( in[52] ) ) - ( $signed( in[94] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_422;
always @( posedge clock ) begin
tree_422 <= ( $signed( in[79] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_423;
always @( posedge clock ) begin
tree_423 <= ( $signed( tree_422 ) ) - ( $signed( tree_61 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_424;
always @( posedge clock ) begin
tree_424 <= ( $signed( in[81] ) ) - ( $signed( in[131] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_425;
always @( posedge clock ) begin
tree_425 <= ( $signed( in[4] ) ) - ( $signed( in[174] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_426;
always @( posedge clock ) begin
tree_426 <= ( $signed( in[76] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_427;
always @( posedge clock ) begin
tree_427 <= ( $signed( tree_426 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_428;
always @( posedge clock ) begin
tree_428 <= ( $signed( tree_427 ) ) - ( $signed( tree_274 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_429;
always @( posedge clock ) begin
tree_429 <= ( $signed( tree_195 ) ) + ( $signed( tree_203 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_430;
always @( posedge clock ) begin
tree_430 <= ( $signed( in[41] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_431;
always @( posedge clock ) begin
tree_431 <= ( $signed( tree_430 ) ) - ( $signed( tree_88 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_432;
always @( posedge clock ) begin
tree_432 <= ( $signed( tree_79 ) ) - ( $signed( tree_64 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_433;
always @( posedge clock ) begin
tree_433 <= ( $signed( tree_30 ) ) + ( $signed( tree_225 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_434;
always @( posedge clock ) begin
tree_434 <= ( $signed( in[21] ) ) - ( $signed( in[142] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_435;
always @( posedge clock ) begin
tree_435 <= ( $signed( in[72] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_436;
always @( posedge clock ) begin
tree_436 <= ( $signed( tree_435 ) ) + ( $signed( tree_187 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_437;
always @( posedge clock ) begin
tree_437 <= ( $signed( in[107] ) ) + ( $signed( in[147] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_438;
always @( posedge clock ) begin
tree_438 <= ( $signed( in[121] ) ) + ( $signed( in[163] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_439;
always @( posedge clock ) begin
tree_439 <= ( $signed( in[42] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_440;
always @( posedge clock ) begin
tree_440 <= ( $signed( tree_439 ) ) + ( $signed( tree_61 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_441;
always @( posedge clock ) begin
tree_441 <= ( $signed( in[8] ) ) - ( $signed( in[80] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_442;
always @( posedge clock ) begin
tree_442 <= ( $signed( in[187] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_443;
always @( posedge clock ) begin
tree_443 <= ( $signed( tree_442 ) ) + ( $signed( tree_37 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_444;
always @( posedge clock ) begin
tree_444 <= ( $signed( tree_5 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_445;
always @( posedge clock ) begin
tree_445 <= ( $signed( tree_444 ) ) + ( $signed( tree_412 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_446;
always @( posedge clock ) begin
tree_446 <= ( $signed( in[70] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_447;
always @( posedge clock ) begin
tree_447 <= ( $signed( tree_446 ) ) - ( $signed( tree_288 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_448;
always @( posedge clock ) begin
tree_448 <= ( $signed( in[125] ) ) - ( $signed( in[130] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_449;
always @( posedge clock ) begin
tree_449 <= ( $signed( in[61] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_450;
always @( posedge clock ) begin
tree_450 <= ( $signed( tree_449 ) ) + ( $signed( tree_176 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_451;
always @( posedge clock ) begin
tree_451 <= ( $signed( in[71] ) ) - ( $signed( in[158] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_452;
always @( posedge clock ) begin
tree_452 <= ( $signed( tree_57 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_453;
always @( posedge clock ) begin
tree_453 <= ( $signed( tree_452 ) ) - ( $signed( tree_410 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_454;
always @( posedge clock ) begin
tree_454 <= ( $signed( in[135] ) ) - ( $signed( in[191] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_455;
always @( posedge clock ) begin
tree_455 <= ( $signed( in[67] ) ) - ( $signed( in[161] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_456;
always @( posedge clock ) begin
tree_456 <= ( $signed( in[40] ) ) + ( $signed( in[124] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_457;
always @( posedge clock ) begin
tree_457 <= ( $signed( tree_408 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_458;
always @( posedge clock ) begin
tree_458 <= ( $signed( tree_457 ) ) + ( $signed( tree_215 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_459;
always @( posedge clock ) begin
tree_459 <= ( $signed( tree_197 ) ) - ( $signed( tree_352 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_460;
always @( posedge clock ) begin
tree_460 <= ( $signed( tree_137 ) ) - ( $signed( tree_382 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_461;
always @( posedge clock ) begin
tree_461 <= ( $signed( in[101] ) ) + ( $signed( in[129] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_462;
always @( posedge clock ) begin
tree_462 <= ( $signed( in[72] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_463;
always @( posedge clock ) begin
tree_463 <= ( $signed( tree_462 ) ) - ( $signed( tree_42 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_464;
always @( posedge clock ) begin
tree_464 <= ( $signed( in[186] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_465;
always @( posedge clock ) begin
tree_465 <= ( $signed( tree_464 ) ) - ( $signed( tree_199 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_466;
always @( posedge clock ) begin
tree_466 <= ( $signed( in[41] ) ) + ( $signed( in[54] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_467;
always @( posedge clock ) begin
tree_467 <= ( $signed( in[57] ) ) - ( $signed( in[142] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_468;
always @( posedge clock ) begin
tree_468 <= ( $signed( tree_19 ) ) + ( $signed( tree_454 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_469;
always @( posedge clock ) begin
tree_469 <= ( $signed( in[3] ) ) - ( $signed( in[187] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_470;
always @( posedge clock ) begin
tree_470 <= ( $signed( in[111] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_471;
always @( posedge clock ) begin
tree_471 <= ( $signed( tree_470 ) ) - ( $signed( tree_152 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_472;
always @( posedge clock ) begin
tree_472 <= ( $signed( tree_79 ) ) - ( $signed( tree_77 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_473;
always @( posedge clock ) begin
tree_473 <= ( $signed( tree_34 ) ) - ( $signed( tree_135 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_474;
always @( posedge clock ) begin
tree_474 <= ( $signed( tree_139 ) ) - ( $signed( tree_6 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_475;
always @( posedge clock ) begin
tree_475 <= ( $signed( in[110] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_476;
always @( posedge clock ) begin
tree_476 <= ( $signed( tree_475 ) ) + ( $signed( tree_145 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_477;
always @( posedge clock ) begin
tree_477 <= ( $signed( in[132] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_478;
always @( posedge clock ) begin
tree_478 <= ( $signed( tree_477 ) ) - ( $signed( tree_62 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_479;
always @( posedge clock ) begin
tree_479 <= ( $signed( tree_87 ) ) + ( $signed( tree_71 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_480;
always @( posedge clock ) begin
tree_480 <= ( $signed( in[68] ) ) - ( $signed( in[72] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_481;
always @( posedge clock ) begin
tree_481 <= ( $signed( in[114] ) ) - ( $signed( in[181] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_482;
always @( posedge clock ) begin
tree_482 <= ( $signed( in[132] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_483;
always @( posedge clock ) begin
tree_483 <= ( $signed( tree_482 ) ) - ( $signed( tree_143 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_484;
always @( posedge clock ) begin
tree_484 <= ( $signed( in[139] ) ) - ( $signed( in[180] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_485;
always @( posedge clock ) begin
tree_485 <= ( $signed( in[21] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_486;
always @( posedge clock ) begin
tree_486 <= ( $signed( tree_485 ) ) - ( $signed( tree_342 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_487;
always @( posedge clock ) begin
tree_487 <= ( $signed( in[9] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_488;
always @( posedge clock ) begin
tree_488 <= ( $signed( tree_487 ) ) - ( $signed( tree_83 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_489;
always @( posedge clock ) begin
tree_489 <= ( $signed( in[23] ) ) - ( $signed( in[43] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_490;
always @( posedge clock ) begin
tree_490 <= ( $signed( in[49] ) ) - ( $signed( in[144] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_491;
always @( posedge clock ) begin
tree_491 <= ( $signed( in[82] ) ) - ( $signed( in[102] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_492;
always @( posedge clock ) begin
tree_492 <= ( $signed( in[55] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_493;
always @( posedge clock ) begin
tree_493 <= ( $signed( tree_492 ) ) - ( $signed( tree_217 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_494;
always @( posedge clock ) begin
tree_494 <= ( $signed( in[139] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_495;
always @( posedge clock ) begin
tree_495 <= ( $signed( tree_494 ) ) - ( $signed( tree_33 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_496;
always @( posedge clock ) begin
tree_496 <= ( $signed( in[6] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_497;
always @( posedge clock ) begin
tree_497 <= ( $signed( tree_496 ) ) + ( $signed( tree_74 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_498;
always @( posedge clock ) begin
tree_498 <= ( $signed( in[54] ) ) - ( $signed( in[65] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_499;
always @( posedge clock ) begin
tree_499 <= ( $signed( in[86] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_500;
always @( posedge clock ) begin
tree_500 <= ( $signed( tree_499 ) ) + ( $signed( tree_1 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_501;
always @( posedge clock ) begin
tree_501 <= ( $signed( in[50] ) ) - ( $signed( in[88] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_502;
always @( posedge clock ) begin
tree_502 <= ( $signed( in[133] ) ) - ( $signed( in[178] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_503;
always @( posedge clock ) begin
tree_503 <= ( $signed( in[16] ) ) + ( $signed( in[59] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_504;
always @( posedge clock ) begin
tree_504 <= ( $signed( tree_192 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_505;
always @( posedge clock ) begin
tree_505 <= ( $signed( tree_504 ) ) + ( $signed( tree_124 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_506;
always @( posedge clock ) begin
tree_506 <= ( $signed( in[61] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_507;
always @( posedge clock ) begin
tree_507 <= ( $signed( tree_506 ) ) - ( $signed( tree_54 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_508;
always @( posedge clock ) begin
tree_508 <= ( $signed( in[116] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_509;
always @( posedge clock ) begin
tree_509 <= ( $signed( tree_508 ) ) - ( $signed( tree_87 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_510;
always @( posedge clock ) begin
tree_510 <= ( $signed( tree_307 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_511;
always @( posedge clock ) begin
tree_511 <=  - ( $signed( tree_510 ) ) + ( $signed( tree_259 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_512;
always @( posedge clock ) begin
tree_512 <= ( $signed( in[164] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_513;
always @( posedge clock ) begin
tree_513 <= ( $signed( tree_512 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_514;
always @( posedge clock ) begin
tree_514 <= ( $signed( tree_513 ) ) + ( $signed( tree_377 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_515;
always @( posedge clock ) begin
tree_515 <= ( $signed( tree_52 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_516;
always @( posedge clock ) begin
tree_516 <= ( $signed( tree_515 ) ) + ( $signed( tree_274 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_517;
always @( posedge clock ) begin
tree_517 <= ( $signed( in[76] ) ) - ( $signed( in[179] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_518;
always @( posedge clock ) begin
tree_518 <= ( $signed( in[31] ) ) - ( $signed( in[81] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_519;
always @( posedge clock ) begin
tree_519 <= ( $signed( in[96] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_520;
always @( posedge clock ) begin
tree_520 <= ( $signed( tree_519 ) ) - ( $signed( tree_75 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_521;
always @( posedge clock ) begin
tree_521 <= ( $signed( in[35] ) ) - ( $signed( in[115] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_522;
always @( posedge clock ) begin
tree_522 <= ( $signed( in[73] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_523;
always @( posedge clock ) begin
tree_523 <= ( $signed( tree_522 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_524;
always @( posedge clock ) begin
tree_524 <= ( $signed( tree_523 ) ) - ( $signed( tree_359 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_525;
always @( posedge clock ) begin
tree_525 <= ( $signed( in[123] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_526;
always @( posedge clock ) begin
tree_526 <= ( $signed( tree_525 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_527;
always @( posedge clock ) begin
tree_527 <= ( $signed( tree_526 ) ) - ( $signed( tree_171 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_528;
always @( posedge clock ) begin
tree_528 <= ( $signed( in[22] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_529;
always @( posedge clock ) begin
tree_529 <= ( $signed( tree_528 ) ) - ( $signed( tree_169 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_530;
always @( posedge clock ) begin
tree_530 <= ( $signed( in[7] ) ) - ( $signed( in[26] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_531;
always @( posedge clock ) begin
tree_531 <= ( $signed( in[122] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_532;
always @( posedge clock ) begin
tree_532 <= ( $signed( tree_531 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_533;
always @( posedge clock ) begin
tree_533 <= ( $signed( tree_532 ) ) - ( $signed( tree_463 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_534;
always @( posedge clock ) begin
tree_534 <= ( $signed( tree_153 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_535;
always @( posedge clock ) begin
tree_535 <= ( $signed( tree_534 ) ) - ( $signed( tree_185 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_536;
always @( posedge clock ) begin
tree_536 <= ( $signed( in[46] ) ) - ( $signed( in[129] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_537;
always @( posedge clock ) begin
tree_537 <= ( $signed( in[127] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_538;
always @( posedge clock ) begin
tree_538 <= ( $signed( tree_537 ) ) - ( $signed( tree_84 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_539;
always @( posedge clock ) begin
tree_539 <= ( $signed( tree_304 ) ) + ( $signed( tree_109 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_540;
always @( posedge clock ) begin
tree_540 <= ( $signed( in[140] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_541;
always @( posedge clock ) begin
tree_541 <= ( $signed( tree_540 ) ) - ( $signed( tree_391 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_542;
always @( posedge clock ) begin
tree_542 <= ( $signed( in[180] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_543;
always @( posedge clock ) begin
tree_543 <= ( $signed( tree_542 ) ) - ( $signed( tree_16 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_544;
always @( posedge clock ) begin
tree_544 <= ( $signed( tree_113 ) ) - ( $signed( tree_281 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_545;
always @( posedge clock ) begin
tree_545 <= ( $signed( in[0] ) ) - ( $signed( in[178] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_546;
always @( posedge clock ) begin
tree_546 <= ( $signed( in[137] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_547;
always @( posedge clock ) begin
tree_547 <= ( $signed( tree_546 ) ) - ( $signed( tree_107 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_548;
always @( posedge clock ) begin
tree_548 <= ( $signed( in[148] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_549;
always @( posedge clock ) begin
tree_549 <= ( $signed( tree_548 ) ) - ( $signed( tree_19 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_550;
always @( posedge clock ) begin
tree_550 <= ( $signed( tree_95 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_551;
always @( posedge clock ) begin
tree_551 <= ( $signed( tree_550 ) ) - ( $signed( tree_282 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_552;
always @( posedge clock ) begin
tree_552 <= ( $signed( in[8] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_553;
always @( posedge clock ) begin
tree_553 <= ( $signed( tree_552 ) ) - ( $signed( tree_32 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_554;
always @( posedge clock ) begin
tree_554 <= ( $signed( in[155] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_555;
always @( posedge clock ) begin
tree_555 <= ( $signed( tree_554 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_556;
always @( posedge clock ) begin
tree_556 <= ( $signed( tree_555 ) ) + ( $signed( tree_340 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_557;
always @( posedge clock ) begin
tree_557 <= ( $signed( in[17] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_558;
always @( posedge clock ) begin
tree_558 <= ( $signed( tree_557 ) ) - ( $signed( tree_60 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_559;
always @( posedge clock ) begin
tree_559 <= ( $signed( in[56] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_560;
always @( posedge clock ) begin
tree_560 <= ( $signed( tree_559 ) ) - ( $signed( tree_138 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_561;
always @( posedge clock ) begin
tree_561 <= ( $signed( in[11] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_562;
always @( posedge clock ) begin
tree_562 <= ( $signed( tree_561 ) ) - ( $signed( tree_244 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_563;
always @( posedge clock ) begin
tree_563 <= ( $signed( in[122] ) ) + ( $signed( in[170] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_564;
always @( posedge clock ) begin
tree_564 <= ( $signed( in[184] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_565;
always @( posedge clock ) begin
tree_565 <= ( $signed( tree_564 ) ) + ( $signed( tree_213 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_566;
always @( posedge clock ) begin
tree_566 <= ( $signed( in[39] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_567;
always @( posedge clock ) begin
tree_567 <= ( $signed( tree_566 ) ) - ( $signed( tree_53 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_568;
always @( posedge clock ) begin
tree_568 <= ( $signed( in[31] ) ) - ( $signed( in[134] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_569;
always @( posedge clock ) begin
tree_569 <= ( $signed( in[48] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_570;
always @( posedge clock ) begin
tree_570 <= ( $signed( tree_569 ) ) - ( $signed( tree_23 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_571;
always @( posedge clock ) begin
tree_571 <= ( $signed( in[71] ) ) - ( $signed( in[190] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_572;
always @( posedge clock ) begin
tree_572 <= ( $signed( tree_71 ) ) - ( $signed( tree_238 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_573;
always @( posedge clock ) begin
tree_573 <= ( $signed( tree_162 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_574;
always @( posedge clock ) begin
tree_574 <= ( $signed( tree_573 ) ) - ( $signed( tree_507 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_575;
always @( posedge clock ) begin
tree_575 <= ( $signed( tree_1 ) ) - ( $signed( tree_298 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_576;
always @( posedge clock ) begin
tree_576 <= ( $signed( tree_52 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_577;
always @( posedge clock ) begin
tree_577 <= ( $signed( tree_576 ) ) - ( $signed( tree_363 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_578;
always @( posedge clock ) begin
tree_578 <= ( $signed( in[32] ) ) - ( $signed( in[87] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_579;
always @( posedge clock ) begin
tree_579 <= ( $signed( tree_330 ) ) + ( $signed( tree_103 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_580;
always @( posedge clock ) begin
tree_580 <= ( $signed( tree_153 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_581;
always @( posedge clock ) begin
tree_581 <= ( $signed( tree_580 ) ) + ( $signed( tree_279 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_582;
always @( posedge clock ) begin
tree_582 <= ( $signed( in[23] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_583;
always @( posedge clock ) begin
tree_583 <= ( $signed( tree_582 ) ) - ( $signed( tree_172 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_584;
always @( posedge clock ) begin
tree_584 <= ( $signed( in[157] ) ) + ( $signed( in[164] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_585;
always @( posedge clock ) begin
tree_585 <= ( $signed( in[26] ) ) - ( $signed( in[183] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_586;
always @( posedge clock ) begin
tree_586 <= ( $signed( in[83] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_587;
always @( posedge clock ) begin
tree_587 <= ( $signed( tree_586 ) ) + ( $signed( tree_131 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_588;
always @( posedge clock ) begin
tree_588 <= ( $signed( in[130] ) ) - ( $signed( in[144] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_589;
always @( posedge clock ) begin
tree_589 <= ( $signed( in[110] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_590;
always @( posedge clock ) begin
tree_590 <= ( $signed( tree_589 ) ) - ( $signed( tree_125 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_591;
always @( posedge clock ) begin
tree_591 <= ( $signed( tree_36 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_592;
always @( posedge clock ) begin
tree_592 <= ( $signed( tree_591 ) ) + ( $signed( tree_556 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_593;
always @( posedge clock ) begin
tree_593 <= ( $signed( in[9] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_594;
always @( posedge clock ) begin
tree_594 <= ( $signed( tree_593 ) ) - ( $signed( tree_28 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_595;
always @( posedge clock ) begin
tree_595 <= ( $signed( in[39] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_596;
always @( posedge clock ) begin
tree_596 <= ( $signed( tree_595 ) ) - ( $signed( tree_341 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_597;
always @( posedge clock ) begin
tree_597 <= ( $signed( in[149] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_598;
always @( posedge clock ) begin
tree_598 <= ( $signed( tree_597 ) ) - ( $signed( tree_327 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_599;
always @( posedge clock ) begin
tree_599 <= ( $signed( in[179] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_600;
always @( posedge clock ) begin
tree_600 <= ( $signed( tree_599 ) ) - ( $signed( tree_568 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_601;
always @( posedge clock ) begin
tree_601 <= ( $signed( in[28] ) ) - ( $signed( in[122] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_602;
always @( posedge clock ) begin
tree_602 <= ( $signed( in[107] ) ) - ( $signed( in[162] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_603;
always @( posedge clock ) begin
tree_603 <= ( $signed( in[42] ) ) - ( $signed( in[95] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_604;
always @( posedge clock ) begin
tree_604 <= ( $signed( in[119] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_605;
always @( posedge clock ) begin
tree_605 <= ( $signed( tree_604 ) ) - ( $signed( tree_95 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_606;
always @( posedge clock ) begin
tree_606 <= ( $signed( in[138] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_607;
always @( posedge clock ) begin
tree_607 <= ( $signed( tree_606 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_608;
always @( posedge clock ) begin
tree_608 <= ( $signed( tree_607 ) ) - ( $signed( tree_465 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_609;
always @( posedge clock ) begin
tree_609 <= ( $signed( in[137] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_610;
always @( posedge clock ) begin
tree_610 <= ( $signed( tree_609 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_611;
always @( posedge clock ) begin
tree_611 <= ( $signed( tree_610 ) ) - ( $signed( tree_479 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_612;
always @( posedge clock ) begin
tree_612 <= ( $signed( tree_38 ) ) - ( $signed( tree_416 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_613;
always @( posedge clock ) begin
tree_613 <= ( $signed( in[64] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_614;
always @( posedge clock ) begin
tree_614 <= ( $signed( tree_613 ) ) - ( $signed( tree_13 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_615;
always @( posedge clock ) begin
tree_615 <= ( $signed( in[117] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_616;
always @( posedge clock ) begin
tree_616 <= ( $signed( tree_615 ) ) - ( $signed( tree_376 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_617;
always @( posedge clock ) begin
tree_617 <= ( $signed( in[18] ) ) + ( $signed( in[111] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_618;
always @( posedge clock ) begin
tree_618 <= ( $signed( in[70] ) ) - ( $signed( in[180] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_619;
always @( posedge clock ) begin
tree_619 <= ( $signed( in[66] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_620;
always @( posedge clock ) begin
tree_620 <= ( $signed( tree_619 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_621;
always @( posedge clock ) begin
tree_621 <= ( $signed( tree_620 ) ) + ( $signed( tree_361 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_622;
always @( posedge clock ) begin
tree_622 <= ( $signed( in[10] ) ) - ( $signed( in[188] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_623;
always @( posedge clock ) begin
tree_623 <= ( $signed( tree_434 ) ) - ( $signed( tree_466 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_624;
always @( posedge clock ) begin
tree_624 <= ( $signed( tree_326 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_625;
always @( posedge clock ) begin
tree_625 <=  - ( $signed( tree_624 ) ) + ( $signed( tree_86 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_626;
always @( posedge clock ) begin
tree_626 <= ( $signed( in[20] ) ) - ( $signed( in[58] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_627;
always @( posedge clock ) begin
tree_627 <= ( $signed( in[48] ) ) - ( $signed( in[97] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_628;
always @( posedge clock ) begin
tree_628 <= ( $signed( in[124] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_629;
always @( posedge clock ) begin
tree_629 <= ( $signed( tree_628 ) ) - ( $signed( tree_115 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_630;
always @( posedge clock ) begin
tree_630 <= ( $signed( in[130] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_631;
always @( posedge clock ) begin
tree_631 <= ( $signed( tree_630 ) ) - ( $signed( tree_289 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_632;
always @( posedge clock ) begin
tree_632 <= ( $signed( in[11] ) ) + ( $signed( in[30] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_633;
always @( posedge clock ) begin
tree_633 <= ( $signed( in[166] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_634;
always @( posedge clock ) begin
tree_634 <= ( $signed( tree_633 ) ) - ( $signed( tree_33 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_635;
always @( posedge clock ) begin
tree_635 <= ( $signed( in[113] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_636;
always @( posedge clock ) begin
tree_636 <= ( $signed( tree_635 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_637;
always @( posedge clock ) begin
tree_637 <= ( $signed( tree_636 ) ) + ( $signed( tree_520 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_638;
always @( posedge clock ) begin
tree_638 <= ( $signed( in[104] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_639;
always @( posedge clock ) begin
tree_639 <= ( $signed( tree_638 ) ) + ( $signed( tree_4 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_640;
always @( posedge clock ) begin
tree_640 <= ( $signed( in[101] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_641;
always @( posedge clock ) begin
tree_641 <= ( $signed( tree_640 ) ) + ( $signed( tree_5 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_642;
always @( posedge clock ) begin
tree_642 <= ( $signed( in[80] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_643;
always @( posedge clock ) begin
tree_643 <= ( $signed( tree_642 ) ) - ( $signed( tree_6 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_644;
always @( posedge clock ) begin
tree_644 <= ( $signed( in[167] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_645;
always @( posedge clock ) begin
tree_645 <= ( $signed( tree_644 ) ) - ( $signed( tree_7 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_646;
always @( posedge clock ) begin
tree_646 <= ( $signed( tree_9 ) ) + ( $signed( tree_10 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_647;
always @( posedge clock ) begin
tree_647 <= ( $signed( tree_11 ) ) + ( $signed( tree_12 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_648;
always @( posedge clock ) begin
tree_648 <= ( $signed( in[28] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_649;
always @( posedge clock ) begin
tree_649 <= ( $signed( tree_648 ) ) - ( $signed( tree_13 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_650;
always @( posedge clock ) begin
tree_650 <= ( $signed( in[50] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_651;
always @( posedge clock ) begin
tree_651 <= ( $signed( tree_650 ) ) - ( $signed( tree_14 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_652;
always @( posedge clock ) begin
tree_652 <= ( $signed( in[99] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_653;
always @( posedge clock ) begin
tree_653 <= ( $signed( tree_652 ) ) - ( $signed( tree_15 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_654;
always @( posedge clock ) begin
tree_654 <= ( $signed( in[185] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_655;
always @( posedge clock ) begin
tree_655 <= ( $signed( tree_654 ) ) - ( $signed( tree_17 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_656;
always @( posedge clock ) begin
tree_656 <= ( $signed( tree_18 ) ) - ( $signed( tree_19 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_657;
always @( posedge clock ) begin
tree_657 <= ( $signed( in[190] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_658;
always @( posedge clock ) begin
tree_658 <= ( $signed( tree_657 ) ) - ( $signed( tree_22 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_659;
always @( posedge clock ) begin
tree_659 <= ( $signed( tree_24 ) ) + ( $signed( tree_25 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_660;
always @( posedge clock ) begin
tree_660 <= ( $signed( in[173] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_661;
always @( posedge clock ) begin
tree_661 <= ( $signed( tree_660 ) ) + ( $signed( tree_26 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_662;
always @( posedge clock ) begin
tree_662 <= ( $signed( in[64] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_663;
always @( posedge clock ) begin
tree_663 <= ( $signed( tree_662 ) ) + ( $signed( tree_27 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_664;
always @( posedge clock ) begin
tree_664 <= ( $signed( in[134] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_665;
always @( posedge clock ) begin
tree_665 <= ( $signed( tree_664 ) ) + ( $signed( tree_28 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_666;
always @( posedge clock ) begin
tree_666 <= ( $signed( in[127] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_667;
always @( posedge clock ) begin
tree_667 <= ( $signed( tree_666 ) ) - ( $signed( tree_29 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_668;
always @( posedge clock ) begin
tree_668 <= ( $signed( in[34] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_669;
always @( posedge clock ) begin
tree_669 <= ( $signed( tree_668 ) ) - ( $signed( tree_30 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_670;
always @( posedge clock ) begin
tree_670 <= ( $signed( in[108] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_671;
always @( posedge clock ) begin
tree_671 <= ( $signed( tree_670 ) ) + ( $signed( tree_34 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_672;
always @( posedge clock ) begin
tree_672 <= ( $signed( tree_28 ) ) + ( $signed( tree_37 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_673;
always @( posedge clock ) begin
tree_673 <= ( $signed( in[91] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_674;
always @( posedge clock ) begin
tree_674 <= ( $signed( tree_673 ) ) - ( $signed( tree_38 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_675;
always @( posedge clock ) begin
tree_675 <= ( $signed( in[181] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_676;
always @( posedge clock ) begin
tree_676 <= ( $signed( tree_675 ) ) + ( $signed( tree_40 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_677;
always @( posedge clock ) begin
tree_677 <= ( $signed( in[57] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_678;
always @( posedge clock ) begin
tree_678 <= ( $signed( tree_677 ) ) - ( $signed( tree_42 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_679;
always @( posedge clock ) begin
tree_679 <= ( $signed( in[115] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_680;
always @( posedge clock ) begin
tree_680 <= ( $signed( tree_679 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_681;
always @( posedge clock ) begin
tree_681 <= ( $signed( tree_680 ) ) - ( $signed( tree_45 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_682;
always @( posedge clock ) begin
tree_682 <= ( $signed( in[179] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_683;
always @( posedge clock ) begin
tree_683 <= ( $signed( tree_682 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_684;
always @( posedge clock ) begin
tree_684 <= ( $signed( tree_683 ) ) - ( $signed( tree_47 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_685;
always @( posedge clock ) begin
tree_685 <= ( $signed( in[172] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_686;
always @( posedge clock ) begin
tree_686 <= ( $signed( tree_685 ) ) - ( $signed( tree_51 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_687;
always @( posedge clock ) begin
tree_687 <= ( $signed( in[94] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_688;
always @( posedge clock ) begin
tree_688 <= ( $signed( tree_687 ) ) + ( $signed( tree_52 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_689;
always @( posedge clock ) begin
tree_689 <= ( $signed( in[22] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_690;
always @( posedge clock ) begin
tree_690 <= ( $signed( tree_689 ) ) - ( $signed( tree_53 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_691;
always @( posedge clock ) begin
tree_691 <= ( $signed( in[12] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_692;
always @( posedge clock ) begin
tree_692 <= ( $signed( tree_691 ) ) - ( $signed( tree_54 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_693;
always @( posedge clock ) begin
tree_693 <= ( $signed( in[42] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_694;
always @( posedge clock ) begin
tree_694 <= ( $signed( tree_693 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_695;
always @( posedge clock ) begin
tree_695 <= ( $signed( tree_694 ) ) + ( $signed( tree_56 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_696;
always @( posedge clock ) begin
tree_696 <= ( $signed( in[29] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_697;
always @( posedge clock ) begin
tree_697 <= ( $signed( tree_696 ) ) - ( $signed( tree_57 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_698;
always @( posedge clock ) begin
tree_698 <= ( $signed( tree_10 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_699;
always @( posedge clock ) begin
tree_699 <= ( $signed( tree_698 ) ) + ( $signed( tree_59 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_700;
always @( posedge clock ) begin
tree_700 <= ( $signed( in[95] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_701;
always @( posedge clock ) begin
tree_701 <= ( $signed( tree_700 ) ) + ( $signed( tree_64 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_702;
always @( posedge clock ) begin
tree_702 <= ( $signed( in[15] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_703;
always @( posedge clock ) begin
tree_703 <= ( $signed( tree_702 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_704;
always @( posedge clock ) begin
tree_704 <= ( $signed( tree_703 ) ) - ( $signed( tree_639 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_705;
always @( posedge clock ) begin
tree_705 <= ( $signed( tree_14 ) ) - ( $signed( tree_65 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_706;
always @( posedge clock ) begin
tree_706 <= ( $signed( in[40] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_707;
always @( posedge clock ) begin
tree_707 <= ( $signed( tree_706 ) ) - ( $signed( tree_71 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_708;
always @( posedge clock ) begin
tree_708 <= ( $signed( in[184] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_709;
always @( posedge clock ) begin
tree_709 <= ( $signed( tree_708 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_710;
always @( posedge clock ) begin
tree_710 <= ( $signed( tree_709 ) ) - ( $signed( tree_73 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_711;
always @( posedge clock ) begin
tree_711 <= ( $signed( in[117] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_712;
always @( posedge clock ) begin
tree_712 <= ( $signed( tree_711 ) ) + ( $signed( tree_75 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_713;
always @( posedge clock ) begin
tree_713 <= ( $signed( in[69] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_714;
always @( posedge clock ) begin
tree_714 <= ( $signed( tree_713 ) ) + ( $signed( tree_76 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_715;
always @( posedge clock ) begin
tree_715 <= ( $signed( tree_78 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_716;
always @( posedge clock ) begin
tree_716 <= ( $signed( tree_715 ) ) + ( $signed( tree_663 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_717;
always @( posedge clock ) begin
tree_717 <= ( $signed( tree_79 ) ) + ( $signed( tree_29 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_718;
always @( posedge clock ) begin
tree_718 <= ( $signed( in[83] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_719;
always @( posedge clock ) begin
tree_719 <= ( $signed( tree_718 ) ) - ( $signed( tree_80 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_720;
always @( posedge clock ) begin
tree_720 <= ( $signed( in[176] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_721;
always @( posedge clock ) begin
tree_721 <= ( $signed( tree_720 ) ) + ( $signed( tree_81 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_722;
always @( posedge clock ) begin
tree_722 <= ( $signed( in[109] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_723;
always @( posedge clock ) begin
tree_723 <= ( $signed( tree_722 ) ) + ( $signed( tree_84 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_724;
always @( posedge clock ) begin
tree_724 <= ( $signed( tree_87 ) ) + ( $signed( tree_88 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_725;
always @( posedge clock ) begin
tree_725 <= ( $signed( tree_75 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_726;
always @( posedge clock ) begin
tree_726 <= ( $signed( tree_725 ) ) + ( $signed( tree_671 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_727;
always @( posedge clock ) begin
tree_727 <= ( $signed( in[58] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_728;
always @( posedge clock ) begin
tree_728 <= ( $signed( tree_727 ) ) - ( $signed( tree_89 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_729;
always @( posedge clock ) begin
tree_729 <= ( $signed( tree_93 ) ) - ( $signed( tree_94 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_730;
always @( posedge clock ) begin
tree_730 <= ( $signed( in[165] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_731;
always @( posedge clock ) begin
tree_731 <= ( $signed( tree_730 ) ) - ( $signed( tree_95 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_732;
always @( posedge clock ) begin
tree_732 <= ( $signed( tree_9 ) ) + ( $signed( tree_96 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_733;
always @( posedge clock ) begin
tree_733 <= ( $signed( in[186] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_734;
always @( posedge clock ) begin
tree_734 <= ( $signed( tree_733 ) ) - ( $signed( tree_97 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_735;
always @( posedge clock ) begin
tree_735 <= ( $signed( tree_639 ) ) - ( $signed( tree_98 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_736;
always @( posedge clock ) begin
tree_736 <= ( $signed( in[47] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_737;
always @( posedge clock ) begin
tree_737 <= ( $signed( tree_736 ) ) - ( $signed( tree_99 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_738;
always @( posedge clock ) begin
tree_738 <= ( $signed( in[78] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_739;
always @( posedge clock ) begin
tree_739 <= ( $signed( tree_738 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_740;
always @( posedge clock ) begin
tree_740 <= ( $signed( tree_739 ) ) + ( $signed( tree_102 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_741;
always @( posedge clock ) begin
tree_741 <= ( $signed( in[5] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_742;
always @( posedge clock ) begin
tree_742 <= ( $signed( tree_741 ) ) - ( $signed( tree_103 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_743;
always @( posedge clock ) begin
tree_743 <= ( $signed( tree_107 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_744;
always @( posedge clock ) begin
tree_744 <=  - ( $signed( tree_743 ) ) + ( $signed( tree_106 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_745;
always @( posedge clock ) begin
tree_745 <= ( $signed( in[63] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_746;
always @( posedge clock ) begin
tree_746 <= ( $signed( tree_745 ) ) - ( $signed( tree_113 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_747;
always @( posedge clock ) begin
tree_747 <= ( $signed( tree_115 ) ) + ( $signed( tree_93 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_748;
always @( posedge clock ) begin
tree_748 <= ( $signed( tree_672 ) ) - ( $signed( tree_117 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_749;
always @( posedge clock ) begin
tree_749 <= ( $signed( tree_118 ) ) - ( $signed( tree_119 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_750;
always @( posedge clock ) begin
tree_750 <= ( $signed( tree_120 ) ) - ( $signed( tree_43 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_751;
always @( posedge clock ) begin
tree_751 <= ( $signed( tree_13 ) ) + ( $signed( tree_121 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_752;
always @( posedge clock ) begin
tree_752 <= ( $signed( in[101] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_753;
always @( posedge clock ) begin
tree_753 <= ( $signed( tree_752 ) ) + ( $signed( tree_122 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_754;
always @( posedge clock ) begin
tree_754 <= ( $signed( tree_53 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_755;
always @( posedge clock ) begin
tree_755 <= ( $signed( tree_754 ) ) - ( $signed( tree_124 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_756;
always @( posedge clock ) begin
tree_756 <= ( $signed( in[143] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_757;
always @( posedge clock ) begin
tree_757 <= ( $signed( tree_756 ) ) - ( $signed( tree_134 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_758;
always @( posedge clock ) begin
tree_758 <= ( $signed( tree_135 ) ) - ( $signed( tree_136 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_759;
always @( posedge clock ) begin
tree_759 <= ( $signed( tree_57 ) ) - ( $signed( tree_137 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_760;
always @( posedge clock ) begin
tree_760 <= ( $signed( tree_60 ) ) - ( $signed( tree_138 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_761;
always @( posedge clock ) begin
tree_761 <= ( $signed( in[92] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_762;
always @( posedge clock ) begin
tree_762 <= ( $signed( tree_761 ) ) - ( $signed( tree_139 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_763;
always @( posedge clock ) begin
tree_763 <= ( $signed( in[21] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_764;
always @( posedge clock ) begin
tree_764 <= ( $signed( tree_763 ) ) + ( $signed( tree_142 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_765;
always @( posedge clock ) begin
tree_765 <= ( $signed( tree_143 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_766;
always @( posedge clock ) begin
tree_766 <= ( $signed( tree_765 ) ) + ( $signed( tree_144 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_767;
always @( posedge clock ) begin
tree_767 <= ( $signed( in[60] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_768;
always @( posedge clock ) begin
tree_768 <= ( $signed( tree_767 ) ) - ( $signed( tree_146 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_769;
always @( posedge clock ) begin
tree_769 <= ( $signed( in[9] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_770;
always @( posedge clock ) begin
tree_770 <= ( $signed( tree_769 ) ) + ( $signed( tree_147 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_771;
always @( posedge clock ) begin
tree_771 <= ( $signed( in[90] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_772;
always @( posedge clock ) begin
tree_772 <= ( $signed( tree_771 ) ) - ( $signed( tree_149 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_773;
always @( posedge clock ) begin
tree_773 <= ( $signed( in[119] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_774;
always @( posedge clock ) begin
tree_774 <= ( $signed( tree_773 ) ) + ( $signed( tree_152 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_775;
always @( posedge clock ) begin
tree_775 <= ( $signed( in[150] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_776;
always @( posedge clock ) begin
tree_776 <= ( $signed( tree_775 ) ) - ( $signed( tree_153 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_777;
always @( posedge clock ) begin
tree_777 <= ( $signed( in[177] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_778;
always @( posedge clock ) begin
tree_778 <= ( $signed( tree_777 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_779;
always @( posedge clock ) begin
tree_779 <= ( $signed( tree_778 ) ) - ( $signed( tree_155 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_780;
always @( posedge clock ) begin
tree_780 <= ( $signed( tree_28 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_781;
always @( posedge clock ) begin
tree_781 <= ( $signed( tree_780 ) ) - ( $signed( tree_159 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_782;
always @( posedge clock ) begin
tree_782 <= ( $signed( in[170] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_783;
always @( posedge clock ) begin
tree_783 <= ( $signed( tree_782 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_784;
always @( posedge clock ) begin
tree_784 <= ( $signed( tree_783 ) ) - ( $signed( tree_731 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_785;
always @( posedge clock ) begin
tree_785 <= ( $signed( in[79] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_786;
always @( posedge clock ) begin
tree_786 <= ( $signed( tree_785 ) ) + ( $signed( tree_161 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_787;
always @( posedge clock ) begin
tree_787 <= ( $signed( in[42] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_788;
always @( posedge clock ) begin
tree_788 <= ( $signed( tree_787 ) ) - ( $signed( tree_162 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_789;
always @( posedge clock ) begin
tree_789 <= ( $signed( in[89] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_790;
always @( posedge clock ) begin
tree_790 <= ( $signed( tree_789 ) ) - ( $signed( tree_163 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_791;
always @( posedge clock ) begin
tree_791 <= ( $signed( tree_165 ) ) + ( $signed( tree_167 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_792;
always @( posedge clock ) begin
tree_792 <= ( $signed( in[95] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_793;
always @( posedge clock ) begin
tree_793 <= ( $signed( tree_792 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_794;
always @( posedge clock ) begin
tree_794 <= ( $signed( tree_793 ) ) - ( $signed( tree_676 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_795;
always @( posedge clock ) begin
tree_795 <= ( $signed( tree_181 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_796;
always @( posedge clock ) begin
tree_796 <= ( $signed( tree_795 ) ) - ( $signed( tree_183 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_797;
always @( posedge clock ) begin
tree_797 <= ( $signed( in[22] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_798;
always @( posedge clock ) begin
tree_798 <= ( $signed( tree_797 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_799;
always @( posedge clock ) begin
tree_799 <= ( $signed( tree_798 ) ) - ( $signed( tree_185 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_800;
always @( posedge clock ) begin
tree_800 <= ( $signed( in[49] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_801;
always @( posedge clock ) begin
tree_801 <= ( $signed( tree_800 ) ) + ( $signed( tree_186 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_802;
always @( posedge clock ) begin
tree_802 <= ( $signed( tree_118 ) ) - ( $signed( tree_191 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_803;
always @( posedge clock ) begin
tree_803 <= ( $signed( in[13] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_804;
always @( posedge clock ) begin
tree_804 <= ( $signed( tree_803 ) ) + ( $signed( tree_195 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_805;
always @( posedge clock ) begin
tree_805 <= ( $signed( in[64] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_806;
always @( posedge clock ) begin
tree_806 <= ( $signed( tree_805 ) ) - ( $signed( tree_196 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_807;
always @( posedge clock ) begin
tree_807 <= ( $signed( in[148] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_808;
always @( posedge clock ) begin
tree_808 <= ( $signed( tree_807 ) ) + ( $signed( tree_197 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_809;
always @( posedge clock ) begin
tree_809 <= ( $signed( tree_15 ) ) - ( $signed( tree_198 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_810;
always @( posedge clock ) begin
tree_810 <= ( $signed( in[58] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_811;
always @( posedge clock ) begin
tree_811 <= ( $signed( tree_810 ) ) + ( $signed( tree_199 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_812;
always @( posedge clock ) begin
tree_812 <= ( $signed( in[93] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_813;
always @( posedge clock ) begin
tree_813 <= ( $signed( tree_812 ) ) - ( $signed( tree_201 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_814;
always @( posedge clock ) begin
tree_814 <= ( $signed( in[191] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_815;
always @( posedge clock ) begin
tree_815 <= ( $signed( tree_814 ) ) - ( $signed( tree_204 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_816;
always @( posedge clock ) begin
tree_816 <= ( $signed( in[106] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_817;
always @( posedge clock ) begin
tree_817 <= ( $signed( tree_816 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_818;
always @( posedge clock ) begin
tree_818 <= ( $signed( tree_817 ) ) + ( $signed( tree_208 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_819;
always @( posedge clock ) begin
tree_819 <= ( $signed( tree_210 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_820;
always @( posedge clock ) begin
tree_820 <= ( $signed( tree_819 ) ) - ( $signed( tree_212 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_821;
always @( posedge clock ) begin
tree_821 <= ( $signed( tree_186 ) ) - ( $signed( tree_213 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_822;
always @( posedge clock ) begin
tree_822 <= ( $signed( tree_216 ) ) - ( $signed( tree_217 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_823;
always @( posedge clock ) begin
tree_823 <= ( $signed( tree_221 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_824;
always @( posedge clock ) begin
tree_824 <= ( $signed( tree_823 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_825;
always @( posedge clock ) begin
tree_825 <= ( $signed( tree_824 ) ) - ( $signed( tree_784 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_826;
always @( posedge clock ) begin
tree_826 <= ( $signed( tree_222 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_827;
always @( posedge clock ) begin
tree_827 <= ( $signed( tree_826 ) ) + ( $signed( tree_224 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_828;
always @( posedge clock ) begin
tree_828 <= ( $signed( tree_146 ) ) - ( $signed( tree_228 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_829;
always @( posedge clock ) begin
tree_829 <= ( $signed( tree_145 ) ) - ( $signed( tree_230 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_830;
always @( posedge clock ) begin
tree_830 <= ( $signed( in[63] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_831;
always @( posedge clock ) begin
tree_831 <= ( $signed( tree_830 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_832;
always @( posedge clock ) begin
tree_832 <= ( $signed( tree_831 ) ) - ( $signed( tree_232 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_833;
always @( posedge clock ) begin
tree_833 <= ( $signed( in[69] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_834;
always @( posedge clock ) begin
tree_834 <= ( $signed( tree_833 ) ) - ( $signed( tree_233 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_835;
always @( posedge clock ) begin
tree_835 <= ( $signed( tree_190 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_836;
always @( posedge clock ) begin
tree_836 <= ( $signed( tree_835 ) ) - ( $signed( tree_237 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_837;
always @( posedge clock ) begin
tree_837 <= ( $signed( tree_7 ) ) - ( $signed( tree_238 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_838;
always @( posedge clock ) begin
tree_838 <= ( $signed( tree_162 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_839;
always @( posedge clock ) begin
tree_839 <= ( $signed( tree_838 ) ) - ( $signed( tree_239 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_840;
always @( posedge clock ) begin
tree_840 <= ( $signed( in[171] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_841;
always @( posedge clock ) begin
tree_841 <= ( $signed( tree_840 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_842;
always @( posedge clock ) begin
tree_842 <= ( $signed( tree_841 ) ) + ( $signed( tree_658 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_843;
always @( posedge clock ) begin
tree_843 <= ( $signed( tree_197 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_844;
always @( posedge clock ) begin
tree_844 <= ( $signed( tree_843 ) ) - ( $signed( tree_774 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_845;
always @( posedge clock ) begin
tree_845 <= ( $signed( in[189] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_846;
always @( posedge clock ) begin
tree_846 <= ( $signed( tree_845 ) ) - ( $signed( tree_254 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_847;
always @( posedge clock ) begin
tree_847 <= ( $signed( tree_89 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_848;
always @( posedge clock ) begin
tree_848 <= ( $signed( tree_847 ) ) - ( $signed( tree_643 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_849;
always @( posedge clock ) begin
tree_849 <= ( $signed( in[100] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_850;
always @( posedge clock ) begin
tree_850 <= ( $signed( tree_849 ) ) + ( $signed( tree_255 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_851;
always @( posedge clock ) begin
tree_851 <= ( $signed( tree_259 ) ) + ( $signed( tree_261 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_852;
always @( posedge clock ) begin
tree_852 <= ( $signed( in[156] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_853;
always @( posedge clock ) begin
tree_853 <= ( $signed( tree_852 ) ) - ( $signed( tree_264 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_854;
always @( posedge clock ) begin
tree_854 <= ( $signed( tree_115 ) ) - ( $signed( tree_265 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_855;
always @( posedge clock ) begin
tree_855 <= ( $signed( tree_94 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_856;
always @( posedge clock ) begin
tree_856 <=  - ( $signed( tree_855 ) ) + ( $signed( tree_274 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_857;
always @( posedge clock ) begin
tree_857 <= ( $signed( in[157] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_858;
always @( posedge clock ) begin
tree_858 <= ( $signed( tree_857 ) ) - ( $signed( tree_276 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_859;
always @( posedge clock ) begin
tree_859 <= ( $signed( tree_277 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_860;
always @( posedge clock ) begin
tree_860 <= ( $signed( tree_859 ) ) + ( $signed( tree_47 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_861;
always @( posedge clock ) begin
tree_861 <= ( $signed( tree_255 ) ) - ( $signed( tree_280 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_862;
always @( posedge clock ) begin
tree_862 <= ( $signed( tree_692 ) ) - ( $signed( tree_285 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_863;
always @( posedge clock ) begin
tree_863 <= ( $signed( in[163] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_864;
always @( posedge clock ) begin
tree_864 <= ( $signed( tree_863 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_865;
always @( posedge clock ) begin
tree_865 <= ( $signed( tree_864 ) ) + ( $signed( tree_672 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_866;
always @( posedge clock ) begin
tree_866 <= ( $signed( in[100] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_867;
always @( posedge clock ) begin
tree_867 <= ( $signed( tree_866 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_868;
always @( posedge clock ) begin
tree_868 <= ( $signed( tree_867 ) ) - ( $signed( tree_639 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_869;
always @( posedge clock ) begin
tree_869 <= ( $signed( in[184] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_870;
always @( posedge clock ) begin
tree_870 <= ( $signed( tree_869 ) ) - ( $signed( tree_298 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_871;
always @( posedge clock ) begin
tree_871 <= ( $signed( tree_301 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_872;
always @( posedge clock ) begin
tree_872 <=  - ( $signed( tree_871 ) ) + ( $signed( tree_663 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_873;
always @( posedge clock ) begin
tree_873 <= ( $signed( tree_200 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_874;
always @( posedge clock ) begin
tree_874 <= ( $signed( tree_873 ) ) + ( $signed( tree_303 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_875;
always @( posedge clock ) begin
tree_875 <= ( $signed( tree_304 ) ) + ( $signed( tree_132 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_876;
always @( posedge clock ) begin
tree_876 <= ( $signed( tree_206 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_877;
always @( posedge clock ) begin
tree_877 <= ( $signed( tree_876 ) ) + ( $signed( tree_306 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_878;
always @( posedge clock ) begin
tree_878 <= ( $signed( in[133] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_879;
always @( posedge clock ) begin
tree_879 <= ( $signed( tree_878 ) ) - ( $signed( tree_316 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_880;
always @( posedge clock ) begin
tree_880 <= ( $signed( tree_319 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_881;
always @( posedge clock ) begin
tree_881 <= ( $signed( tree_880 ) ) - ( $signed( tree_321 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_882;
always @( posedge clock ) begin
tree_882 <= ( $signed( in[18] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_883;
always @( posedge clock ) begin
tree_883 <= ( $signed( tree_882 ) ) + ( $signed( tree_322 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_884;
always @( posedge clock ) begin
tree_884 <= ( $signed( tree_324 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_885;
always @( posedge clock ) begin
tree_885 <= ( $signed( tree_884 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_886;
always @( posedge clock ) begin
tree_886 <= ( $signed( tree_885 ) ) - ( $signed( tree_249 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_887;
always @( posedge clock ) begin
tree_887 <= ( $signed( tree_330 ) ) + ( $signed( tree_331 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_888;
always @( posedge clock ) begin
tree_888 <= ( $signed( in[83] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_889;
always @( posedge clock ) begin
tree_889 <= ( $signed( tree_888 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_890;
always @( posedge clock ) begin
tree_890 <= ( $signed( tree_889 ) ) - ( $signed( tree_336 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_891;
always @( posedge clock ) begin
tree_891 <= ( $signed( tree_168 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_892;
always @( posedge clock ) begin
tree_892 <= ( $signed( tree_891 ) ) - ( $signed( tree_815 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_893;
always @( posedge clock ) begin
tree_893 <= ( $signed( tree_307 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_894;
always @( posedge clock ) begin
tree_894 <= ( $signed( tree_893 ) ) + ( $signed( tree_340 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_895;
always @( posedge clock ) begin
tree_895 <= ( $signed( in[43] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_896;
always @( posedge clock ) begin
tree_896 <= ( $signed( tree_895 ) ) - ( $signed( tree_343 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_897;
always @( posedge clock ) begin
tree_897 <= ( $signed( tree_352 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_898;
always @( posedge clock ) begin
tree_898 <= ( $signed( tree_897 ) ) - ( $signed( tree_354 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_899;
always @( posedge clock ) begin
tree_899 <= ( $signed( tree_357 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_900;
always @( posedge clock ) begin
tree_900 <=  - ( $signed( tree_899 ) ) + ( $signed( tree_356 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_901;
always @( posedge clock ) begin
tree_901 <= ( $signed( in[15] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_902;
always @( posedge clock ) begin
tree_902 <= ( $signed( tree_901 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_903;
always @( posedge clock ) begin
tree_903 <= ( $signed( tree_902 ) ) + ( $signed( tree_645 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_904;
always @( posedge clock ) begin
tree_904 <= ( $signed( tree_216 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_905;
always @( posedge clock ) begin
tree_905 <= ( $signed( tree_904 ) ) + ( $signed( tree_728 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_906;
always @( posedge clock ) begin
tree_906 <= ( $signed( tree_4 ) ) - ( $signed( tree_358 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_907;
always @( posedge clock ) begin
tree_907 <= ( $signed( in[39] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_908;
always @( posedge clock ) begin
tree_908 <= ( $signed( tree_907 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_909;
always @( posedge clock ) begin
tree_909 <= ( $signed( tree_908 ) ) - ( $signed( tree_690 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_910;
always @( posedge clock ) begin
tree_910 <= ( $signed( in[14] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_911;
always @( posedge clock ) begin
tree_911 <= ( $signed( tree_910 ) ) - ( $signed( tree_365 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_912;
always @( posedge clock ) begin
tree_912 <= ( $signed( tree_213 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_913;
always @( posedge clock ) begin
tree_913 <= ( $signed( tree_912 ) ) + ( $signed( tree_639 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_914;
always @( posedge clock ) begin
tree_914 <= ( $signed( tree_135 ) ) + ( $signed( tree_374 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_915;
always @( posedge clock ) begin
tree_915 <= ( $signed( tree_724 ) ) + ( $signed( tree_375 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_916;
always @( posedge clock ) begin
tree_916 <= ( $signed( in[82] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_917;
always @( posedge clock ) begin
tree_917 <= ( $signed( tree_916 ) ) - ( $signed( tree_382 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_918;
always @( posedge clock ) begin
tree_918 <= ( $signed( in[180] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_919;
always @( posedge clock ) begin
tree_919 <= ( $signed( tree_918 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_920;
always @( posedge clock ) begin
tree_920 <= ( $signed( tree_919 ) ) - ( $signed( tree_712 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_921;
always @( posedge clock ) begin
tree_921 <= ( $signed( in[110] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_922;
always @( posedge clock ) begin
tree_922 <= ( $signed( tree_921 ) ) + ( $signed( tree_387 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_923;
always @( posedge clock ) begin
tree_923 <= ( $signed( tree_330 ) ) + ( $signed( tree_388 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_924;
always @( posedge clock ) begin
tree_924 <= ( $signed( tree_99 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_925;
always @( posedge clock ) begin
tree_925 <= ( $signed( tree_924 ) ) - ( $signed( tree_397 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_926;
always @( posedge clock ) begin
tree_926 <= ( $signed( in[89] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_927;
always @( posedge clock ) begin
tree_927 <= ( $signed( tree_926 ) ) + ( $signed( tree_398 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_928;
always @( posedge clock ) begin
tree_928 <= ( $signed( tree_319 ) ) + ( $signed( tree_403 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_929;
always @( posedge clock ) begin
tree_929 <= ( $signed( tree_404 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_930;
always @( posedge clock ) begin
tree_930 <= ( $signed( tree_929 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_931;
always @( posedge clock ) begin
tree_931 <= ( $signed( tree_930 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_932;
always @( posedge clock ) begin
tree_932 <= ( $signed( tree_931 ) ) - ( $signed( tree_407 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_933;
always @( posedge clock ) begin
tree_933 <= ( $signed( tree_669 ) ) - ( $signed( tree_98 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_934;
always @( posedge clock ) begin
tree_934 <= ( $signed( tree_308 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_935;
always @( posedge clock ) begin
tree_935 <=  - ( $signed( tree_934 ) ) + ( $signed( tree_412 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_936;
always @( posedge clock ) begin
tree_936 <= ( $signed( tree_63 ) ) - ( $signed( tree_416 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_937;
always @( posedge clock ) begin
tree_937 <= ( $signed( in[168] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_938;
always @( posedge clock ) begin
tree_938 <= ( $signed( tree_937 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_939;
always @( posedge clock ) begin
tree_939 <= ( $signed( tree_938 ) ) + ( $signed( tree_418 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_940;
always @( posedge clock ) begin
tree_940 <= ( $signed( in[175] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_941;
always @( posedge clock ) begin
tree_941 <= ( $signed( tree_940 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_942;
always @( posedge clock ) begin
tree_942 <= ( $signed( tree_941 ) ) - ( $signed( tree_712 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_943;
always @( posedge clock ) begin
tree_943 <= ( $signed( tree_191 ) ) - ( $signed( tree_425 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_944;
always @( posedge clock ) begin
tree_944 <= ( $signed( tree_139 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_945;
always @( posedge clock ) begin
tree_945 <= ( $signed( tree_944 ) ) - ( $signed( tree_645 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_946;
always @( posedge clock ) begin
tree_946 <= ( $signed( tree_434 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_947;
always @( posedge clock ) begin
tree_947 <= ( $signed( tree_946 ) ) + ( $signed( tree_436 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_948;
always @( posedge clock ) begin
tree_948 <= ( $signed( in[133] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_949;
always @( posedge clock ) begin
tree_949 <= ( $signed( tree_948 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_950;
always @( posedge clock ) begin
tree_950 <= ( $signed( tree_949 ) ) - ( $signed( tree_788 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_951;
always @( posedge clock ) begin
tree_951 <= ( $signed( tree_714 ) ) + ( $signed( tree_359 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_952;
always @( posedge clock ) begin
tree_952 <= ( $signed( tree_438 ) ) - ( $signed( tree_316 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_953;
always @( posedge clock ) begin
tree_953 <= ( $signed( in[55] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_954;
always @( posedge clock ) begin
tree_954 <= ( $signed( tree_953 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_955;
always @( posedge clock ) begin
tree_955 <= ( $signed( tree_954 ) ) + ( $signed( tree_443 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_956;
always @( posedge clock ) begin
tree_956 <= ( $signed( tree_175 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_957;
always @( posedge clock ) begin
tree_957 <= ( $signed( tree_956 ) ) + ( $signed( tree_447 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_958;
always @( posedge clock ) begin
tree_958 <= ( $signed( in[188] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_959;
always @( posedge clock ) begin
tree_959 <= ( $signed( tree_958 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_960;
always @( posedge clock ) begin
tree_960 <= ( $signed( tree_959 ) ) + ( $signed( tree_717 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_961;
always @( posedge clock ) begin
tree_961 <= ( $signed( in[90] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_962;
always @( posedge clock ) begin
tree_962 <= ( $signed( tree_961 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_963;
always @( posedge clock ) begin
tree_963 <= ( $signed( tree_962 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_964;
always @( posedge clock ) begin
tree_964 <= ( $signed( tree_963 ) ) - ( $signed( tree_920 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_965;
always @( posedge clock ) begin
tree_965 <= ( $signed( in[129] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_966;
always @( posedge clock ) begin
tree_966 <= ( $signed( tree_965 ) ) - ( $signed( tree_448 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_967;
always @( posedge clock ) begin
tree_967 <= ( $signed( tree_24 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_968;
always @( posedge clock ) begin
tree_968 <= ( $signed( tree_967 ) ) + ( $signed( tree_641 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_969;
always @( posedge clock ) begin
tree_969 <= ( $signed( tree_195 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_970;
always @( posedge clock ) begin
tree_970 <= ( $signed( tree_969 ) ) + ( $signed( tree_721 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_971;
always @( posedge clock ) begin
tree_971 <= ( $signed( in[170] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_972;
always @( posedge clock ) begin
tree_972 <= ( $signed( tree_971 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_973;
always @( posedge clock ) begin
tree_973 <= ( $signed( tree_972 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_974;
always @( posedge clock ) begin
tree_974 <= ( $signed( tree_973 ) ) - ( $signed( tree_681 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_975;
always @( posedge clock ) begin
tree_975 <= ( $signed( tree_451 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_976;
always @( posedge clock ) begin
tree_976 <= ( $signed( tree_975 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_977;
always @( posedge clock ) begin
tree_977 <= ( $signed( tree_976 ) ) + ( $signed( tree_453 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_978;
always @( posedge clock ) begin
tree_978 <= ( $signed( tree_6 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_979;
always @( posedge clock ) begin
tree_979 <= ( $signed( tree_978 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_980;
always @( posedge clock ) begin
tree_980 <= ( $signed( tree_979 ) ) - ( $signed( tree_458 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_981;
always @( posedge clock ) begin
tree_981 <= ( $signed( tree_461 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_982;
always @( posedge clock ) begin
tree_982 <=  - ( $signed( tree_981 ) ) + ( $signed( tree_321 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_983;
always @( posedge clock ) begin
tree_983 <= ( $signed( tree_655 ) ) - ( $signed( tree_379 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_984;
always @( posedge clock ) begin
tree_984 <= ( $signed( in[36] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_985;
always @( posedge clock ) begin
tree_985 <= ( $signed( tree_984 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_986;
always @( posedge clock ) begin
tree_986 <= ( $signed( tree_985 ) ) + ( $signed( tree_674 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_987;
always @( posedge clock ) begin
tree_987 <= ( $signed( tree_658 ) ) - ( $signed( tree_697 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_988;
always @( posedge clock ) begin
tree_988 <= ( $signed( tree_438 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_989;
always @( posedge clock ) begin
tree_989 <= ( $signed( tree_988 ) ) + ( $signed( tree_478 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_990;
always @( posedge clock ) begin
tree_990 <= ( $signed( in[45] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_991;
always @( posedge clock ) begin
tree_991 <= ( $signed( tree_990 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_992;
always @( posedge clock ) begin
tree_992 <= ( $signed( tree_991 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_993;
always @( posedge clock ) begin
tree_993 <= ( $signed( tree_992 ) ) - ( $signed( tree_726 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_994;
always @( posedge clock ) begin
tree_994 <= ( $signed( tree_17 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_995;
always @( posedge clock ) begin
tree_995 <= ( $signed( tree_994 ) ) - ( $signed( tree_483 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_996;
always @( posedge clock ) begin
tree_996 <= ( $signed( tree_448 ) ) - ( $signed( tree_484 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_997;
always @( posedge clock ) begin
tree_997 <= ( $signed( in[97] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_998;
always @( posedge clock ) begin
tree_998 <= ( $signed( tree_997 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_999;
always @( posedge clock ) begin
tree_999 <= ( $signed( tree_998 ) ) + ( $signed( tree_486 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1000;
always @( posedge clock ) begin
tree_1000 <= ( $signed( in[145] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1001;
always @( posedge clock ) begin
tree_1001 <= ( $signed( tree_1000 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1002;
always @( posedge clock ) begin
tree_1002 <= ( $signed( tree_1001 ) ) + ( $signed( tree_896 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1003;
always @( posedge clock ) begin
tree_1003 <= ( $signed( tree_246 ) ) + ( $signed( tree_488 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1004;
always @( posedge clock ) begin
tree_1004 <= ( $signed( tree_714 ) ) - ( $signed( tree_768 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1005;
always @( posedge clock ) begin
tree_1005 <= ( $signed( tree_490 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1006;
always @( posedge clock ) begin
tree_1006 <= ( $signed( tree_1005 ) ) - ( $signed( tree_440 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1007;
always @( posedge clock ) begin
tree_1007 <= ( $signed( in[151] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1008;
always @( posedge clock ) begin
tree_1008 <= ( $signed( tree_1007 ) ) + ( $signed( tree_491 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1009;
always @( posedge clock ) begin
tree_1009 <= ( $signed( tree_327 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1010;
always @( posedge clock ) begin
tree_1010 <=  - ( $signed( tree_1009 ) ) + ( $signed( tree_731 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1011;
always @( posedge clock ) begin
tree_1011 <= ( $signed( in[162] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1012;
always @( posedge clock ) begin
tree_1012 <= ( $signed( tree_1011 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1013;
always @( posedge clock ) begin
tree_1013 <= ( $signed( tree_1012 ) ) + ( $signed( tree_500 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1014;
always @( posedge clock ) begin
tree_1014 <= ( $signed( tree_328 ) ) - ( $signed( tree_502 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1015;
always @( posedge clock ) begin
tree_1015 <= ( $signed( in[40] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1016;
always @( posedge clock ) begin
tree_1016 <= ( $signed( tree_1015 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1017;
always @( posedge clock ) begin
tree_1017 <= ( $signed( tree_1016 ) ) + ( $signed( tree_770 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1018;
always @( posedge clock ) begin
tree_1018 <= ( $signed( tree_420 ) ) + ( $signed( tree_659 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1019;
always @( posedge clock ) begin
tree_1019 <= ( $signed( tree_172 ) ) + ( $signed( tree_517 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1020;
always @( posedge clock ) begin
tree_1020 <= ( $signed( tree_104 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1021;
always @( posedge clock ) begin
tree_1021 <= ( $signed( tree_1020 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1022;
always @( posedge clock ) begin
tree_1022 <= ( $signed( tree_1021 ) ) - ( $signed( tree_524 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1023;
always @( posedge clock ) begin
tree_1023 <= ( $signed( tree_529 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1024;
always @( posedge clock ) begin
tree_1024 <=  - ( $signed( tree_1023 ) ) + ( $signed( tree_527 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1025;
always @( posedge clock ) begin
tree_1025 <= ( $signed( tree_54 ) ) + ( $signed( tree_530 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1026;
always @( posedge clock ) begin
tree_1026 <= ( $signed( in[155] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1027;
always @( posedge clock ) begin
tree_1027 <= ( $signed( tree_1026 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1028;
always @( posedge clock ) begin
tree_1028 <= ( $signed( tree_1027 ) ) - ( $signed( tree_669 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1029;
always @( posedge clock ) begin
tree_1029 <= ( $signed( in[12] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1030;
always @( posedge clock ) begin
tree_1030 <= ( $signed( tree_1029 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1031;
always @( posedge clock ) begin
tree_1031 <= ( $signed( tree_1030 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1032;
always @( posedge clock ) begin
tree_1032 <= ( $signed( tree_1031 ) ) - ( $signed( tree_535 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1033;
always @( posedge clock ) begin
tree_1033 <= ( $signed( tree_22 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1034;
always @( posedge clock ) begin
tree_1034 <= ( $signed( tree_1033 ) ) - ( $signed( tree_538 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1035;
always @( posedge clock ) begin
tree_1035 <= ( $signed( tree_544 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1036;
always @( posedge clock ) begin
tree_1036 <=  - ( $signed( tree_1035 ) ) + ( $signed( tree_960 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1037;
always @( posedge clock ) begin
tree_1037 <= ( $signed( tree_465 ) ) - ( $signed( tree_553 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1038;
always @( posedge clock ) begin
tree_1038 <= ( $signed( in[125] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1039;
always @( posedge clock ) begin
tree_1039 <= ( $signed( tree_1038 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1040;
always @( posedge clock ) begin
tree_1040 <= ( $signed( tree_1039 ) ) + ( $signed( tree_562 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1041;
always @( posedge clock ) begin
tree_1041 <= ( $signed( tree_565 ) ) + ( $signed( tree_567 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1042;
always @( posedge clock ) begin
tree_1042 <= ( $signed( tree_377 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1043;
always @( posedge clock ) begin
tree_1043 <= ( $signed( tree_1042 ) ) - ( $signed( tree_577 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1044;
always @( posedge clock ) begin
tree_1044 <= ( $signed( tree_578 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1045;
always @( posedge clock ) begin
tree_1045 <= ( $signed( tree_1044 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1046;
always @( posedge clock ) begin
tree_1046 <= ( $signed( tree_1045 ) ) - ( $signed( tree_935 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1047;
always @( posedge clock ) begin
tree_1047 <= ( $signed( tree_37 ) ) - ( $signed( tree_584 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1048;
always @( posedge clock ) begin
tree_1048 <= ( $signed( tree_585 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1049;
always @( posedge clock ) begin
tree_1049 <=  - ( $signed( tree_1048 ) ) + ( $signed( tree_707 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1050;
always @( posedge clock ) begin
tree_1050 <= ( $signed( in[136] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1051;
always @( posedge clock ) begin
tree_1051 <= ( $signed( tree_1050 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1052;
always @( posedge clock ) begin
tree_1052 <= ( $signed( tree_1051 ) ) - ( $signed( tree_887 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1053;
always @( posedge clock ) begin
tree_1053 <= ( $signed( tree_590 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1054;
always @( posedge clock ) begin
tree_1054 <=  - ( $signed( tree_1053 ) ) + ( $signed( tree_842 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1055;
always @( posedge clock ) begin
tree_1055 <= ( $signed( tree_280 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1056;
always @( posedge clock ) begin
tree_1056 <= ( $signed( tree_1055 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1057;
always @( posedge clock ) begin
tree_1057 <= ( $signed( tree_1056 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1058;
always @( posedge clock ) begin
tree_1058 <= ( $signed( tree_1057 ) ) + ( $signed( tree_592 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1059;
always @( posedge clock ) begin
tree_1059 <= ( $signed( tree_0 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1060;
always @( posedge clock ) begin
tree_1060 <= ( $signed( tree_1059 ) ) - ( $signed( tree_714 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1061;
always @( posedge clock ) begin
tree_1061 <= ( $signed( tree_495 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1062;
always @( posedge clock ) begin
tree_1062 <= ( $signed( tree_1061 ) ) + ( $signed( tree_621 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1063;
always @( posedge clock ) begin
tree_1063 <= ( $signed( in[4] ) ) + ( $signed( in[36] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1064;
always @( posedge clock ) begin
tree_1064 <= ( $signed( in[95] ) ) + ( $signed( in[130] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1065;
always @( posedge clock ) begin
tree_1065 <= ( $signed( tree_1063 ) ) + ( $signed( tree_1064 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1066;
always @( posedge clock ) begin
tree_1066 <= ( $signed( tree_146 ) ) - ( $signed( tree_136 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1067;
always @( posedge clock ) begin
tree_1067 <= ( $signed( tree_403 ) ) - ( $signed( tree_181 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1068;
always @( posedge clock ) begin
tree_1068 <= ( $signed( tree_617 ) ) + ( $signed( tree_456 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1069;
always @( posedge clock ) begin
tree_1069 <= ( $signed( tree_1065 ) ) + ( $signed( tree_1066 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1070;
always @( posedge clock ) begin
tree_1070 <= ( $signed( tree_1067 ) ) + ( $signed( tree_1068 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1071;
always @( posedge clock ) begin
tree_1071 <=  - ( $signed( tree_447 ) ) + ( $signed( tree_861 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1072;
always @( posedge clock ) begin
tree_1072 <= ( $signed( tree_688 ) ) + ( $signed( tree_560 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1073;
always @( posedge clock ) begin
tree_1073 <= ( $signed( tree_1069 ) ) + ( $signed( tree_1070 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1074;
always @( posedge clock ) begin
tree_1074 <= ( $signed( tree_1071 ) ) + ( $signed( tree_1072 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1075;
always @( posedge clock ) begin
tree_1075 <= ( $signed( tree_842 ) ) + ( $signed( tree_868 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1076;
always @( posedge clock ) begin
tree_1076 <= ( $signed( tree_1052 ) ) + ( $signed( tree_925 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1077;
always @( posedge clock ) begin
tree_1077 <= ( $signed( tree_955 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1078;
always @( posedge clock ) begin
tree_1078 <= ( $signed( tree_1073 ) ) + ( $signed( tree_1074 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1079;
always @( posedge clock ) begin
tree_1079 <= ( $signed( tree_1075 ) ) + ( $signed( tree_1076 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1080;
always @( posedge clock ) begin
tree_1080 <= ( $signed( tree_1077 ) ) + ( $signed( tree_1032 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1081;
always @( posedge clock ) begin
tree_1081 <= ( $signed( tree_1062 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1082;
always @( posedge clock ) begin
tree_1082 <= ( $signed( tree_1078 ) ) + ( $signed( tree_1079 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1083;
always @( posedge clock ) begin
tree_1083 <= ( $signed( tree_1080 ) ) + ( $signed( tree_1081 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1084;
always @( posedge clock ) begin
tree_1084 <= ( $signed( tree_1082 ) ) + ( $signed( tree_1083 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1085;
always @( posedge clock ) begin
tree_1085 <= ( $signed( tree_622 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1086;
always @( posedge clock ) begin
tree_1086 <= ( $signed( tree_1085 ) ) - ( $signed( tree_623 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1087;
always @( posedge clock ) begin
tree_1087 <= ( $signed( tree_269 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1088;
always @( posedge clock ) begin
tree_1088 <= ( $signed( tree_1087 ) ) + ( $signed( tree_625 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1089;
always @( posedge clock ) begin
tree_1089 <= ( $signed( tree_632 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1090;
always @( posedge clock ) begin
tree_1090 <= ( $signed( tree_1089 ) ) - ( $signed( tree_634 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1091;
always @( posedge clock ) begin
tree_1091 <= ( $signed( in[0] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1092;
always @( posedge clock ) begin
tree_1092 <= ( $signed( tree_1091 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1093;
always @( posedge clock ) begin
tree_1093 <= ( $signed( tree_1092 ) ) + ( $signed( tree_639 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1094;
always @( posedge clock ) begin
tree_1094 <= ( $signed( in[163] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1095;
always @( posedge clock ) begin
tree_1095 <= ( $signed( tree_1094 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1096;
always @( posedge clock ) begin
tree_1096 <= ( $signed( tree_1095 ) ) - ( $signed( tree_645 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1097;
always @( posedge clock ) begin
tree_1097 <= ( $signed( tree_16 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1098;
always @( posedge clock ) begin
tree_1098 <= ( $signed( tree_1097 ) ) - ( $signed( tree_655 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1099;
always @( posedge clock ) begin
tree_1099 <= ( $signed( tree_21 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1100;
always @( posedge clock ) begin
tree_1100 <= ( $signed( tree_1099 ) ) - ( $signed( tree_658 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1101;
always @( posedge clock ) begin
tree_1101 <= ( $signed( tree_23 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1102;
always @( posedge clock ) begin
tree_1102 <= ( $signed( tree_1101 ) ) - ( $signed( tree_659 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1103;
always @( posedge clock ) begin
tree_1103 <= ( $signed( tree_663 ) ) + ( $signed( tree_665 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1104;
always @( posedge clock ) begin
tree_1104 <= ( $signed( tree_31 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1105;
always @( posedge clock ) begin
tree_1105 <=  - ( $signed( tree_1104 ) ) + ( $signed( tree_669 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1106;
always @( posedge clock ) begin
tree_1106 <= ( $signed( in[138] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1107;
always @( posedge clock ) begin
tree_1107 <= ( $signed( tree_1106 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1108;
always @( posedge clock ) begin
tree_1108 <= ( $signed( tree_1107 ) ) + ( $signed( tree_672 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1109;
always @( posedge clock ) begin
tree_1109 <= ( $signed( tree_41 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1110;
always @( posedge clock ) begin
tree_1110 <= ( $signed( tree_1109 ) ) + ( $signed( tree_678 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1111;
always @( posedge clock ) begin
tree_1111 <= ( $signed( tree_690 ) ) - ( $signed( tree_692 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1112;
always @( posedge clock ) begin
tree_1112 <= ( $signed( in[5] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1113;
always @( posedge clock ) begin
tree_1113 <= ( $signed( tree_1112 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1114;
always @( posedge clock ) begin
tree_1114 <= ( $signed( tree_1113 ) ) - ( $signed( tree_697 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1115;
always @( posedge clock ) begin
tree_1115 <= ( $signed( tree_63 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1116;
always @( posedge clock ) begin
tree_1116 <= ( $signed( tree_1115 ) ) + ( $signed( tree_701 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1117;
always @( posedge clock ) begin
tree_1117 <= ( $signed( in[160] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1118;
always @( posedge clock ) begin
tree_1118 <= ( $signed( tree_1117 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1119;
always @( posedge clock ) begin
tree_1119 <= ( $signed( tree_1118 ) ) - ( $signed( tree_705 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1120;
always @( posedge clock ) begin
tree_1120 <= ( $signed( in[161] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1121;
always @( posedge clock ) begin
tree_1121 <= ( $signed( tree_1120 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1122;
always @( posedge clock ) begin
tree_1122 <= ( $signed( tree_1121 ) ) - ( $signed( tree_707 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1123;
always @( posedge clock ) begin
tree_1123 <= ( $signed( in[115] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1124;
always @( posedge clock ) begin
tree_1124 <= ( $signed( tree_1123 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1125;
always @( posedge clock ) begin
tree_1125 <= ( $signed( tree_1124 ) ) + ( $signed( tree_712 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1126;
always @( posedge clock ) begin
tree_1126 <= ( $signed( tree_18 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1127;
always @( posedge clock ) begin
tree_1127 <= ( $signed( tree_1126 ) ) - ( $signed( tree_714 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1128;
always @( posedge clock ) begin
tree_1128 <= ( $signed( tree_77 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1129;
always @( posedge clock ) begin
tree_1129 <= ( $signed( tree_1128 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1130;
always @( posedge clock ) begin
tree_1130 <= ( $signed( tree_1129 ) ) - ( $signed( tree_716 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1131;
always @( posedge clock ) begin
tree_1131 <= ( $signed( in[138] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1132;
always @( posedge clock ) begin
tree_1132 <= ( $signed( tree_1131 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1133;
always @( posedge clock ) begin
tree_1133 <= ( $signed( tree_1132 ) ) - ( $signed( tree_717 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1134;
always @( posedge clock ) begin
tree_1134 <= ( $signed( in[71] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1135;
always @( posedge clock ) begin
tree_1135 <= ( $signed( tree_1134 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1136;
always @( posedge clock ) begin
tree_1136 <= ( $signed( tree_1135 ) ) + ( $signed( tree_721 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1137;
always @( posedge clock ) begin
tree_1137 <= ( $signed( tree_83 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1138;
always @( posedge clock ) begin
tree_1138 <= ( $signed( tree_1137 ) ) + ( $signed( tree_723 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1139;
always @( posedge clock ) begin
tree_1139 <= ( $signed( tree_2 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1140;
always @( posedge clock ) begin
tree_1140 <= ( $signed( tree_1139 ) ) - ( $signed( tree_724 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1141;
always @( posedge clock ) begin
tree_1141 <= ( $signed( tree_731 ) ) + ( $signed( tree_732 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1142;
always @( posedge clock ) begin
tree_1142 <= ( $signed( tree_45 ) ) - ( $signed( tree_737 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1143;
always @( posedge clock ) begin
tree_1143 <= ( $signed( tree_5 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1144;
always @( posedge clock ) begin
tree_1144 <= ( $signed( tree_1143 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1145;
always @( posedge clock ) begin
tree_1145 <= ( $signed( tree_1144 ) ) + ( $signed( tree_740 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1146;
always @( posedge clock ) begin
tree_1146 <= ( $signed( tree_104 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1147;
always @( posedge clock ) begin
tree_1147 <= ( $signed( tree_1146 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1148;
always @( posedge clock ) begin
tree_1148 <= ( $signed( tree_1147 ) ) - ( $signed( tree_744 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1149;
always @( posedge clock ) begin
tree_1149 <= ( $signed( in[102] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1150;
always @( posedge clock ) begin
tree_1150 <= ( $signed( tree_1149 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1151;
always @( posedge clock ) begin
tree_1151 <= ( $signed( tree_1150 ) ) - ( $signed( tree_747 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1152;
always @( posedge clock ) begin
tree_1152 <= ( $signed( tree_753 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1153;
always @( posedge clock ) begin
tree_1153 <= ( $signed( tree_1152 ) ) + ( $signed( tree_755 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1154;
always @( posedge clock ) begin
tree_1154 <= ( $signed( tree_78 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1155;
always @( posedge clock ) begin
tree_1155 <= ( $signed( tree_1154 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1156;
always @( posedge clock ) begin
tree_1156 <= ( $signed( tree_1155 ) ) - ( $signed( tree_1125 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1157;
always @( posedge clock ) begin
tree_1157 <= ( $signed( in[144] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1158;
always @( posedge clock ) begin
tree_1158 <= ( $signed( tree_1157 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1159;
always @( posedge clock ) begin
tree_1159 <= ( $signed( tree_1158 ) ) - ( $signed( tree_758 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1160;
always @( posedge clock ) begin
tree_1160 <= ( $signed( tree_65 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1161;
always @( posedge clock ) begin
tree_1161 <= ( $signed( tree_1160 ) ) - ( $signed( tree_759 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1162;
always @( posedge clock ) begin
tree_1162 <= ( $signed( tree_762 ) ) - ( $signed( tree_141 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1163;
always @( posedge clock ) begin
tree_1163 <= ( $signed( in[2] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1164;
always @( posedge clock ) begin
tree_1164 <= ( $signed( tree_1163 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1165;
always @( posedge clock ) begin
tree_1165 <= ( $signed( tree_1164 ) ) + ( $signed( tree_770 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1166;
always @( posedge clock ) begin
tree_1166 <= ( $signed( in[131] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1167;
always @( posedge clock ) begin
tree_1167 <= ( $signed( tree_1166 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1168;
always @( posedge clock ) begin
tree_1168 <= ( $signed( tree_1167 ) ) - ( $signed( tree_774 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1169;
always @( posedge clock ) begin
tree_1169 <= ( $signed( in[152] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1170;
always @( posedge clock ) begin
tree_1170 <= ( $signed( tree_1169 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1171;
always @( posedge clock ) begin
tree_1171 <= ( $signed( tree_1170 ) ) - ( $signed( tree_776 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1172;
always @( posedge clock ) begin
tree_1172 <= ( $signed( tree_83 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1173;
always @( posedge clock ) begin
tree_1173 <= ( $signed( tree_1172 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1174;
always @( posedge clock ) begin
tree_1174 <= ( $signed( tree_1173 ) ) - ( $signed( tree_784 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1175;
always @( posedge clock ) begin
tree_1175 <= ( $signed( in[141] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1176;
always @( posedge clock ) begin
tree_1176 <= ( $signed( tree_1175 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1177;
always @( posedge clock ) begin
tree_1177 <= ( $signed( tree_1176 ) ) + ( $signed( tree_788 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1178;
always @( posedge clock ) begin
tree_1178 <= ( $signed( tree_641 ) ) + ( $signed( tree_790 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1179;
always @( posedge clock ) begin
tree_1179 <= ( $signed( in[179] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1180;
always @( posedge clock ) begin
tree_1180 <= ( $signed( tree_1179 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1181;
always @( posedge clock ) begin
tree_1181 <= ( $signed( tree_1180 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1182;
always @( posedge clock ) begin
tree_1182 <= ( $signed( tree_1181 ) ) + ( $signed( tree_799 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1183;
always @( posedge clock ) begin
tree_1183 <= ( $signed( tree_165 ) ) + ( $signed( tree_801 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1184;
always @( posedge clock ) begin
tree_1184 <= ( $signed( in[101] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1185;
always @( posedge clock ) begin
tree_1185 <= ( $signed( tree_1184 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1186;
always @( posedge clock ) begin
tree_1186 <= ( $signed( tree_1185 ) ) - ( $signed( tree_808 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1187;
always @( posedge clock ) begin
tree_1187 <= ( $signed( tree_200 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1188;
always @( posedge clock ) begin
tree_1188 <= ( $signed( tree_1187 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1189;
always @( posedge clock ) begin
tree_1189 <=  - ( $signed( tree_1188 ) ) + ( $signed( tree_1093 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1190;
always @( posedge clock ) begin
tree_1190 <= ( $signed( tree_3 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1191;
always @( posedge clock ) begin
tree_1191 <= ( $signed( tree_1190 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1192;
always @( posedge clock ) begin
tree_1192 <= ( $signed( tree_1191 ) ) + ( $signed( tree_1108 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1193;
always @( posedge clock ) begin
tree_1193 <= ( $signed( tree_215 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1194;
always @( posedge clock ) begin
tree_1194 <=  - ( $signed( tree_1193 ) ) + ( $signed( tree_1093 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1195;
always @( posedge clock ) begin
tree_1195 <= ( $signed( tree_220 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1196;
always @( posedge clock ) begin
tree_1196 <= ( $signed( tree_1195 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1197;
always @( posedge clock ) begin
tree_1197 <= ( $signed( tree_1196 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1198;
always @( posedge clock ) begin
tree_1198 <= ( $signed( tree_1197 ) ) - ( $signed( tree_825 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1199;
always @( posedge clock ) begin
tree_1199 <= ( $signed( tree_828 ) ) - ( $signed( tree_802 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1200;
always @( posedge clock ) begin
tree_1200 <= ( $signed( in[40] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1201;
always @( posedge clock ) begin
tree_1201 <= ( $signed( tree_1200 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1202;
always @( posedge clock ) begin
tree_1202 <= ( $signed( tree_1201 ) ) - ( $signed( tree_829 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1203;
always @( posedge clock ) begin
tree_1203 <= ( $signed( in[165] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1204;
always @( posedge clock ) begin
tree_1204 <= ( $signed( tree_1203 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1205;
always @( posedge clock ) begin
tree_1205 <= ( $signed( tree_1204 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1206;
always @( posedge clock ) begin
tree_1206 <= ( $signed( tree_1205 ) ) - ( $signed( tree_836 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1207;
always @( posedge clock ) begin
tree_1207 <= ( $signed( tree_240 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1208;
always @( posedge clock ) begin
tree_1208 <= ( $signed( tree_1207 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1209;
always @( posedge clock ) begin
tree_1209 <= ( $signed( tree_1208 ) ) - ( $signed( tree_1156 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1210;
always @( posedge clock ) begin
tree_1210 <= ( $signed( in[27] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1211;
always @( posedge clock ) begin
tree_1211 <= ( $signed( tree_1210 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1212;
always @( posedge clock ) begin
tree_1212 <= ( $signed( tree_1211 ) ) + ( $signed( tree_850 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1213;
always @( posedge clock ) begin
tree_1213 <= ( $signed( tree_257 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1214;
always @( posedge clock ) begin
tree_1214 <= ( $signed( tree_1213 ) ) + ( $signed( tree_851 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1215;
always @( posedge clock ) begin
tree_1215 <= ( $signed( tree_853 ) ) - ( $signed( tree_854 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1216;
always @( posedge clock ) begin
tree_1216 <= ( $signed( tree_275 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1217;
always @( posedge clock ) begin
tree_1217 <= ( $signed( tree_1216 ) ) - ( $signed( tree_858 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1218;
always @( posedge clock ) begin
tree_1218 <= ( $signed( in[164] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1219;
always @( posedge clock ) begin
tree_1219 <= ( $signed( tree_1218 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1220;
always @( posedge clock ) begin
tree_1220 <= ( $signed( tree_1219 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1221;
always @( posedge clock ) begin
tree_1221 <= ( $signed( tree_1220 ) ) - ( $signed( tree_1096 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1222;
always @( posedge clock ) begin
tree_1222 <= ( $signed( tree_287 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1223;
always @( posedge clock ) begin
tree_1223 <=  - ( $signed( tree_1222 ) ) + ( $signed( tree_865 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1224;
always @( posedge clock ) begin
tree_1224 <= ( $signed( in[1] ) ) + ( $signed( in[24] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1225;
always @( posedge clock ) begin
tree_1225 <=  - ( $signed( in[89] ) ) + ( $signed( in[138] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1226;
always @( posedge clock ) begin
tree_1226 <= ( $signed( in[141] ) ) + ( $signed( in[146] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1227;
always @( posedge clock ) begin
tree_1227 <= ( $signed( in[181] ) ) + ( $signed( in[185] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1228;
always @( posedge clock ) begin
tree_1228 <= ( $signed( tree_1224 ) ) + ( $signed( tree_1225 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1229;
always @( posedge clock ) begin
tree_1229 <= ( $signed( tree_1226 ) ) + ( $signed( tree_1227 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1230;
always @( posedge clock ) begin
tree_1230 <=  - ( $signed( tree_37 ) ) + ( $signed( tree_139 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1231;
always @( posedge clock ) begin
tree_1231 <= ( $signed( tree_199 ) ) + ( $signed( tree_216 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1232;
always @( posedge clock ) begin
tree_1232 <=  - ( $signed( tree_288 ) ) + ( $signed( tree_265 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1233;
always @( posedge clock ) begin
tree_1233 <=  - ( $signed( tree_289 ) ) + ( $signed( tree_51 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1234;
always @( posedge clock ) begin
tree_1234 <= ( $signed( tree_131 ) ) - ( $signed( tree_293 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1235;
always @( posedge clock ) begin
tree_1235 <= ( $signed( tree_296 ) ) + ( $signed( tree_297 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1236;
always @( posedge clock ) begin
tree_1236 <= ( $signed( tree_1228 ) ) - ( $signed( tree_1229 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1237;
always @( posedge clock ) begin
tree_1237 <= ( $signed( tree_1230 ) ) + ( $signed( tree_1231 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1238;
always @( posedge clock ) begin
tree_1238 <= ( $signed( tree_1232 ) ) + ( $signed( tree_1233 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1239;
always @( posedge clock ) begin
tree_1239 <= ( $signed( tree_1234 ) ) - ( $signed( tree_1235 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1240;
always @( posedge clock ) begin
tree_1240 <= ( $signed( tree_701 ) ) + ( $signed( tree_240 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1241;
always @( posedge clock ) begin
tree_1241 <= ( $signed( tree_861 ) ) + ( $signed( tree_808 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1242;
always @( posedge clock ) begin
tree_1242 <= ( $signed( tree_295 ) ) - ( $signed( tree_870 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1243;
always @( posedge clock ) begin
tree_1243 <= ( $signed( tree_875 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1244;
always @( posedge clock ) begin
tree_1244 <= ( $signed( tree_1236 ) ) + ( $signed( tree_1237 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1245;
always @( posedge clock ) begin
tree_1245 <= ( $signed( tree_1238 ) ) + ( $signed( tree_1239 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1246;
always @( posedge clock ) begin
tree_1246 <=  - ( $signed( tree_1240 ) ) + ( $signed( tree_1241 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1247;
always @( posedge clock ) begin
tree_1247 <= ( $signed( tree_1242 ) ) + ( $signed( tree_1243 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1248;
always @( posedge clock ) begin
tree_1248 <= ( $signed( tree_292 ) ) + ( $signed( tree_868 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1249;
always @( posedge clock ) begin
tree_1249 <=  - ( $signed( tree_300 ) ) + ( $signed( tree_872 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1250;
always @( posedge clock ) begin
tree_1250 <=  - ( $signed( tree_874 ) ) + ( $signed( tree_877 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1251;
always @( posedge clock ) begin
tree_1251 <= ( $signed( tree_1244 ) ) + ( $signed( tree_1245 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1252;
always @( posedge clock ) begin
tree_1252 <= ( $signed( tree_1246 ) ) + ( $signed( tree_1247 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1253;
always @( posedge clock ) begin
tree_1253 <=  - ( $signed( tree_1248 ) ) + ( $signed( tree_1249 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1254;
always @( posedge clock ) begin
tree_1254 <= ( $signed( tree_1250 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1255;
always @( posedge clock ) begin
tree_1255 <= ( $signed( tree_1251 ) ) + ( $signed( tree_1252 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1256;
always @( posedge clock ) begin
tree_1256 <= ( $signed( tree_1253 ) ) + ( $signed( tree_1254 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1257;
always @( posedge clock ) begin
tree_1257 <= ( $signed( tree_1255 ) ) + ( $signed( tree_1256 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1258;
always @( posedge clock ) begin
tree_1258 <= ( $signed( in[141] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1259;
always @( posedge clock ) begin
tree_1259 <= ( $signed( tree_1258 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1260;
always @( posedge clock ) begin
tree_1260 <= ( $signed( tree_1259 ) ) - ( $signed( tree_883 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1261;
always @( posedge clock ) begin
tree_1261 <= ( $signed( tree_671 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1262;
always @( posedge clock ) begin
tree_1262 <= ( $signed( tree_1261 ) ) + ( $signed( tree_894 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1263;
always @( posedge clock ) begin
tree_1263 <= ( $signed( tree_205 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1264;
always @( posedge clock ) begin
tree_1264 <= ( $signed( tree_1263 ) ) + ( $signed( tree_906 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1265;
always @( posedge clock ) begin
tree_1265 <= ( $signed( tree_232 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1266;
always @( posedge clock ) begin
tree_1266 <= ( $signed( tree_1265 ) ) - ( $signed( tree_1116 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1267;
always @( posedge clock ) begin
tree_1267 <= ( $signed( in[32] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1268;
always @( posedge clock ) begin
tree_1268 <= ( $signed( tree_1267 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1269;
always @( posedge clock ) begin
tree_1269 <= ( $signed( tree_1268 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1270;
always @( posedge clock ) begin
tree_1270 <= ( $signed( tree_1269 ) ) + ( $signed( tree_920 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1271;
always @( posedge clock ) begin
tree_1271 <= ( $signed( tree_390 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1272;
always @( posedge clock ) begin
tree_1272 <= ( $signed( tree_1271 ) ) + ( $signed( tree_1140 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1273;
always @( posedge clock ) begin
tree_1273 <= ( $signed( tree_244 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1274;
always @( posedge clock ) begin
tree_1274 <= ( $signed( tree_1273 ) ) - ( $signed( tree_927 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1275;
always @( posedge clock ) begin
tree_1275 <= ( $signed( tree_401 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1276;
always @( posedge clock ) begin
tree_1276 <=  - ( $signed( tree_1275 ) ) + ( $signed( tree_1199 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1277;
always @( posedge clock ) begin
tree_1277 <= ( $signed( tree_818 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1278;
always @( posedge clock ) begin
tree_1278 <= ( $signed( tree_1277 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1279;
always @( posedge clock ) begin
tree_1279 <= ( $signed( tree_1278 ) ) + ( $signed( tree_932 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1280;
always @( posedge clock ) begin
tree_1280 <= ( $signed( tree_96 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1281;
always @( posedge clock ) begin
tree_1281 <= ( $signed( tree_1280 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1282;
always @( posedge clock ) begin
tree_1282 <= ( $signed( tree_1281 ) ) + ( $signed( tree_942 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1283;
always @( posedge clock ) begin
tree_1283 <= ( $signed( tree_933 ) ) - ( $signed( tree_945 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1284;
always @( posedge clock ) begin
tree_1284 <= ( $signed( tree_433 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1285;
always @( posedge clock ) begin
tree_1285 <=  - ( $signed( tree_1284 ) ) + ( $signed( tree_1093 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1286;
always @( posedge clock ) begin
tree_1286 <= ( $signed( in[4] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1287;
always @( posedge clock ) begin
tree_1287 <= ( $signed( tree_1286 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1288;
always @( posedge clock ) begin
tree_1288 <= ( $signed( tree_1287 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1289;
always @( posedge clock ) begin
tree_1289 <= ( $signed( tree_1288 ) ) + ( $signed( tree_947 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1290;
always @( posedge clock ) begin
tree_1290 <= ( $signed( tree_129 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1291;
always @( posedge clock ) begin
tree_1291 <= ( $signed( tree_1290 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1292;
always @( posedge clock ) begin
tree_1292 <= ( $signed( tree_1291 ) ) + ( $signed( tree_950 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1293;
always @( posedge clock ) begin
tree_1293 <= ( $signed( tree_1110 ) ) + ( $signed( tree_951 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1294;
always @( posedge clock ) begin
tree_1294 <= ( $signed( tree_329 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1295;
always @( posedge clock ) begin
tree_1295 <= ( $signed( tree_1294 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1296;
always @( posedge clock ) begin
tree_1296 <= ( $signed( tree_1295 ) ) + ( $signed( tree_957 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1297;
always @( posedge clock ) begin
tree_1297 <= ( $signed( in[92] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1298;
always @( posedge clock ) begin
tree_1298 <= ( $signed( tree_1297 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1299;
always @( posedge clock ) begin
tree_1299 <= ( $signed( tree_1298 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1300;
always @( posedge clock ) begin
tree_1300 <= ( $signed( tree_1299 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1301;
always @( posedge clock ) begin
tree_1301 <= ( $signed( tree_1300 ) ) - ( $signed( tree_964 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1302;
always @( posedge clock ) begin
tree_1302 <= ( $signed( in[19] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1303;
always @( posedge clock ) begin
tree_1303 <= ( $signed( tree_1302 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1304;
always @( posedge clock ) begin
tree_1304 <= ( $signed( tree_1303 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1305;
always @( posedge clock ) begin
tree_1305 <= ( $signed( tree_1304 ) ) + ( $signed( tree_968 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1306;
always @( posedge clock ) begin
tree_1306 <= ( $signed( tree_142 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1307;
always @( posedge clock ) begin
tree_1307 <= ( $signed( tree_1306 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1308;
always @( posedge clock ) begin
tree_1308 <= ( $signed( tree_1307 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1309;
always @( posedge clock ) begin
tree_1309 <= ( $signed( tree_1308 ) ) + ( $signed( tree_974 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1310;
always @( posedge clock ) begin
tree_1310 <= ( $signed( in[153] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1311;
always @( posedge clock ) begin
tree_1311 <= ( $signed( tree_1310 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1312;
always @( posedge clock ) begin
tree_1312 <= ( $signed( tree_1311 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1313;
always @( posedge clock ) begin
tree_1313 <= ( $signed( tree_1312 ) ) + ( $signed( tree_1125 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1314;
always @( posedge clock ) begin
tree_1314 <= ( $signed( in[10] ) ) + ( $signed( in[62] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1315;
always @( posedge clock ) begin
tree_1315 <= ( $signed( in[75] ) ) + ( $signed( in[81] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1316;
always @( posedge clock ) begin
tree_1316 <= ( $signed( in[166] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1317;
always @( posedge clock ) begin
tree_1317 <=  - ( $signed( tree_1314 ) ) + ( $signed( tree_1315 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1318;
always @( posedge clock ) begin
tree_1318 <= ( $signed( tree_1316 ) ) + ( $signed( tree_22 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1319;
always @( posedge clock ) begin
tree_1319 <= ( $signed( tree_20 ) ) - ( $signed( tree_15 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1320;
always @( posedge clock ) begin
tree_1320 <= ( $signed( tree_213 ) ) + ( $signed( tree_288 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1321;
always @( posedge clock ) begin
tree_1321 <= ( $signed( tree_466 ) ) - ( $signed( tree_480 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1322;
always @( posedge clock ) begin
tree_1322 <= ( $signed( tree_481 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1323;
always @( posedge clock ) begin
tree_1323 <= ( $signed( tree_1317 ) ) - ( $signed( tree_1318 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1324;
always @( posedge clock ) begin
tree_1324 <= ( $signed( tree_1319 ) ) - ( $signed( tree_1320 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1325;
always @( posedge clock ) begin
tree_1325 <= ( $signed( tree_1321 ) ) - ( $signed( tree_1322 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1326;
always @( posedge clock ) begin
tree_1326 <=  - ( $signed( tree_336 ) ) + ( $signed( tree_345 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1327;
always @( posedge clock ) begin
tree_1327 <= ( $signed( tree_479 ) ) - ( $signed( tree_996 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1328;
always @( posedge clock ) begin
tree_1328 <= ( $signed( tree_750 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1329;
always @( posedge clock ) begin
tree_1329 <= ( $signed( tree_1323 ) ) + ( $signed( tree_1324 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1330;
always @( posedge clock ) begin
tree_1330 <= ( $signed( tree_1325 ) ) + ( $signed( tree_1326 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1331;
always @( posedge clock ) begin
tree_1331 <= ( $signed( tree_1327 ) ) - ( $signed( tree_1328 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1332;
always @( posedge clock ) begin
tree_1332 <= ( $signed( tree_844 ) ) + ( $signed( tree_995 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1333;
always @( posedge clock ) begin
tree_1333 <=  - ( $signed( tree_999 ) ) + ( $signed( tree_1002 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1334;
always @( posedge clock ) begin
tree_1334 <= ( $signed( tree_1003 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1335;
always @( posedge clock ) begin
tree_1335 <= ( $signed( tree_1329 ) ) + ( $signed( tree_1330 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1336;
always @( posedge clock ) begin
tree_1336 <= ( $signed( tree_1331 ) ) - ( $signed( tree_1332 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1337;
always @( posedge clock ) begin
tree_1337 <= ( $signed( tree_1333 ) ) - ( $signed( tree_1334 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1338;
always @( posedge clock ) begin
tree_1338 <= ( $signed( tree_993 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1339;
always @( posedge clock ) begin
tree_1339 <= ( $signed( tree_1335 ) ) + ( $signed( tree_1336 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1340;
always @( posedge clock ) begin
tree_1340 <= ( $signed( tree_1337 ) ) - ( $signed( tree_1338 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1341;
always @( posedge clock ) begin
tree_1341 <= ( $signed( tree_1339 ) ) + ( $signed( tree_1340 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1342;
always @( posedge clock ) begin
tree_1342 <= ( $signed( in[31] ) ) + ( $signed( in[37] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1343;
always @( posedge clock ) begin
tree_1343 <= ( $signed( in[49] ) ) + ( $signed( in[100] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1344;
always @( posedge clock ) begin
tree_1344 <= ( $signed( in[176] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1345;
always @( posedge clock ) begin
tree_1345 <= ( $signed( tree_1342 ) ) + ( $signed( tree_1343 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1346;
always @( posedge clock ) begin
tree_1346 <= ( $signed( tree_1344 ) ) - ( $signed( tree_197 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1347;
always @( posedge clock ) begin
tree_1347 <= ( $signed( tree_204 ) ) + ( $signed( tree_358 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1348;
always @( posedge clock ) begin
tree_1348 <= ( $signed( tree_227 ) ) - ( $signed( tree_413 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1349;
always @( posedge clock ) begin
tree_1349 <= ( $signed( tree_498 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1350;
always @( posedge clock ) begin
tree_1350 <= ( $signed( tree_1345 ) ) + ( $signed( tree_1346 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1351;
always @( posedge clock ) begin
tree_1351 <= ( $signed( tree_1347 ) ) + ( $signed( tree_1348 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1352;
always @( posedge clock ) begin
tree_1352 <= ( $signed( tree_1349 ) ) + ( $signed( tree_641 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1353;
always @( posedge clock ) begin
tree_1353 <=  - ( $signed( tree_412 ) ) + ( $signed( tree_732 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1354;
always @( posedge clock ) begin
tree_1354 <=  - ( $signed( tree_433 ) ) + ( $signed( tree_493 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1355;
always @( posedge clock ) begin
tree_1355 <= ( $signed( tree_495 ) ) - ( $signed( tree_497 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1356;
always @( posedge clock ) begin
tree_1356 <= ( $signed( tree_1350 ) ) + ( $signed( tree_1351 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1357;
always @( posedge clock ) begin
tree_1357 <=  - ( $signed( tree_1352 ) ) + ( $signed( tree_1353 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1358;
always @( posedge clock ) begin
tree_1358 <= ( $signed( tree_1354 ) ) + ( $signed( tree_1355 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1359;
always @( posedge clock ) begin
tree_1359 <= ( $signed( tree_704 ) ) + ( $signed( tree_947 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1360;
always @( posedge clock ) begin
tree_1360 <= ( $signed( tree_839 ) ) - ( $signed( tree_1010 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1361;
always @( posedge clock ) begin
tree_1361 <= ( $signed( tree_862 ) ) + ( $signed( tree_1013 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1362;
always @( posedge clock ) begin
tree_1362 <= ( $signed( tree_1356 ) ) + ( $signed( tree_1357 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1363;
always @( posedge clock ) begin
tree_1363 <= ( $signed( tree_1358 ) ) + ( $signed( tree_1359 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1364;
always @( posedge clock ) begin
tree_1364 <= ( $signed( tree_1360 ) ) + ( $signed( tree_1361 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1365;
always @( posedge clock ) begin
tree_1365 <= ( $signed( tree_1362 ) ) + ( $signed( tree_1363 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1366;
always @( posedge clock ) begin
tree_1366 <= ( $signed( tree_1364 ) ) + ( $signed( tree_1301 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1367;
always @( posedge clock ) begin
tree_1367 <= ( $signed( tree_1365 ) ) + ( $signed( tree_1366 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1368;
always @( posedge clock ) begin
tree_1368 <= ( $signed( in[51] ) ) + ( $signed( in[84] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1369;
always @( posedge clock ) begin
tree_1369 <= ( $signed( in[117] ) ) - ( $signed( in[165] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1370;
always @( posedge clock ) begin
tree_1370 <=  - ( $signed( tree_1368 ) ) + ( $signed( tree_1369 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1371;
always @( posedge clock ) begin
tree_1371 <= ( $signed( tree_38 ) ) + ( $signed( tree_195 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1372;
always @( posedge clock ) begin
tree_1372 <= ( $signed( tree_1 ) ) - ( $signed( tree_230 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1373;
always @( posedge clock ) begin
tree_1373 <= ( $signed( tree_324 ) ) + ( $signed( tree_501 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1374;
always @( posedge clock ) begin
tree_1374 <= ( $signed( tree_503 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1375;
always @( posedge clock ) begin
tree_1375 <= ( $signed( tree_1370 ) ) - ( $signed( tree_1371 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1376;
always @( posedge clock ) begin
tree_1376 <= ( $signed( tree_1372 ) ) + ( $signed( tree_1373 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1377;
always @( posedge clock ) begin
tree_1377 <=  - ( $signed( tree_1374 ) ) + ( $signed( tree_714 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1378;
always @( posedge clock ) begin
tree_1378 <= ( $signed( tree_47 ) ) + ( $signed( tree_212 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1379;
always @( posedge clock ) begin
tree_1379 <=  - ( $signed( tree_381 ) ) + ( $signed( tree_373 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1380;
always @( posedge clock ) begin
tree_1380 <= ( $signed( tree_1014 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1381;
always @( posedge clock ) begin
tree_1381 <= ( $signed( tree_1375 ) ) + ( $signed( tree_1376 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1382;
always @( posedge clock ) begin
tree_1382 <= ( $signed( tree_1377 ) ) + ( $signed( tree_1378 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1383;
always @( posedge clock ) begin
tree_1383 <= ( $signed( tree_1379 ) ) - ( $signed( tree_1380 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1384;
always @( posedge clock ) begin
tree_1384 <= ( $signed( tree_844 ) ) + ( $signed( tree_796 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1385;
always @( posedge clock ) begin
tree_1385 <= ( $signed( tree_1017 ) ) + ( $signed( tree_905 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1386;
always @( posedge clock ) begin
tree_1386 <= ( $signed( tree_505 ) ) + ( $signed( tree_1018 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1387;
always @( posedge clock ) begin
tree_1387 <= ( $signed( tree_1381 ) ) + ( $signed( tree_1382 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1388;
always @( posedge clock ) begin
tree_1388 <= ( $signed( tree_1383 ) ) - ( $signed( tree_1384 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1389;
always @( posedge clock ) begin
tree_1389 <= ( $signed( tree_1385 ) ) + ( $signed( tree_1386 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1390;
always @( posedge clock ) begin
tree_1390 <= ( $signed( tree_1387 ) ) + ( $signed( tree_1388 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1391;
always @( posedge clock ) begin
tree_1391 <= ( $signed( tree_1389 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1392;
always @( posedge clock ) begin
tree_1392 <= ( $signed( tree_1390 ) ) - ( $signed( tree_1391 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1393;
always @( posedge clock ) begin
tree_1393 <= ( $signed( in[38] ) ) + ( $signed( in[78] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1394;
always @( posedge clock ) begin
tree_1394 <= ( $signed( in[147] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1395;
always @( posedge clock ) begin
tree_1395 <= ( $signed( tree_1393 ) ) + ( $signed( tree_1394 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1396;
always @( posedge clock ) begin
tree_1396 <=  - ( $signed( tree_27 ) ) + ( $signed( tree_19 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1397;
always @( posedge clock ) begin
tree_1397 <= ( $signed( tree_38 ) ) + ( $signed( tree_42 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1398;
always @( posedge clock ) begin
tree_1398 <= ( $signed( tree_118 ) ) + ( $signed( tree_15 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1399;
always @( posedge clock ) begin
tree_1399 <= ( $signed( tree_341 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1400;
always @( posedge clock ) begin
tree_1400 <= ( $signed( tree_1395 ) ) + ( $signed( tree_1396 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1401;
always @( posedge clock ) begin
tree_1401 <= ( $signed( tree_1397 ) ) - ( $signed( tree_1398 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1402;
always @( posedge clock ) begin
tree_1402 <=  - ( $signed( tree_1399 ) ) + ( $signed( tree_507 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1403;
always @( posedge clock ) begin
tree_1403 <=  - ( $signed( tree_311 ) ) + ( $signed( tree_429 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1404;
always @( posedge clock ) begin
tree_1404 <=  - ( $signed( tree_509 ) ) + ( $signed( tree_996 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1405;
always @( posedge clock ) begin
tree_1405 <= ( $signed( tree_1019 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1406;
always @( posedge clock ) begin
tree_1406 <= ( $signed( tree_1400 ) ) + ( $signed( tree_1401 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1407;
always @( posedge clock ) begin
tree_1407 <= ( $signed( tree_1402 ) ) + ( $signed( tree_1403 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1408;
always @( posedge clock ) begin
tree_1408 <= ( $signed( tree_1404 ) ) + ( $signed( tree_1405 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1409;
always @( posedge clock ) begin
tree_1409 <=  - ( $signed( tree_511 ) ) + ( $signed( tree_514 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1410;
always @( posedge clock ) begin
tree_1410 <= ( $signed( tree_516 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1411;
always @( posedge clock ) begin
tree_1411 <= ( $signed( tree_1406 ) ) + ( $signed( tree_1407 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1412;
always @( posedge clock ) begin
tree_1412 <= ( $signed( tree_1408 ) ) + ( $signed( tree_1409 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1413;
always @( posedge clock ) begin
tree_1413 <= ( $signed( tree_1410 ) ) + ( $signed( tree_1283 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1414;
always @( posedge clock ) begin
tree_1414 <= ( $signed( tree_1411 ) ) + ( $signed( tree_1412 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1415;
always @( posedge clock ) begin
tree_1415 <= ( $signed( tree_1413 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1416;
always @( posedge clock ) begin
tree_1416 <= ( $signed( tree_1414 ) ) + ( $signed( tree_1415 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1417;
always @( posedge clock ) begin
tree_1417 <= ( $signed( in[32] ) ) + ( $signed( in[34] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1418;
always @( posedge clock ) begin
tree_1418 <= ( $signed( in[52] ) ) + ( $signed( in[108] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1419;
always @( posedge clock ) begin
tree_1419 <= ( $signed( in[161] ) ) - ( $signed( in[189] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1420;
always @( posedge clock ) begin
tree_1420 <= ( $signed( tree_1417 ) ) + ( $signed( tree_1418 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1421;
always @( posedge clock ) begin
tree_1421 <= ( $signed( tree_1419 ) ) - ( $signed( tree_152 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1422;
always @( posedge clock ) begin
tree_1422 <= ( $signed( tree_200 ) ) + ( $signed( tree_196 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1423;
always @( posedge clock ) begin
tree_1423 <= ( $signed( tree_518 ) ) + ( $signed( tree_521 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1424;
always @( posedge clock ) begin
tree_1424 <= ( $signed( tree_48 ) ) + ( $signed( tree_325 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1425;
always @( posedge clock ) begin
tree_1425 <=  - ( $signed( tree_1420 ) ) + ( $signed( tree_1421 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1426;
always @( posedge clock ) begin
tree_1426 <=  - ( $signed( tree_1422 ) ) + ( $signed( tree_1423 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1427;
always @( posedge clock ) begin
tree_1427 <= ( $signed( tree_1424 ) ) + ( $signed( tree_185 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1428;
always @( posedge clock ) begin
tree_1428 <= ( $signed( tree_285 ) ) + ( $signed( tree_758 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1429;
always @( posedge clock ) begin
tree_1429 <= ( $signed( tree_659 ) ) - ( $signed( tree_167 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1430;
always @( posedge clock ) begin
tree_1430 <=  - ( $signed( tree_345 ) ) + ( $signed( tree_520 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1431;
always @( posedge clock ) begin
tree_1431 <= ( $signed( tree_180 ) ) - ( $signed( tree_1025 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1432;
always @( posedge clock ) begin
tree_1432 <= ( $signed( tree_1425 ) ) + ( $signed( tree_1426 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1433;
always @( posedge clock ) begin
tree_1433 <= ( $signed( tree_1427 ) ) + ( $signed( tree_1428 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1434;
always @( posedge clock ) begin
tree_1434 <= ( $signed( tree_1429 ) ) + ( $signed( tree_1430 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1435;
always @( posedge clock ) begin
tree_1435 <= ( $signed( tree_1431 ) ) + ( $signed( tree_1127 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1436;
always @( posedge clock ) begin
tree_1436 <= ( $signed( tree_1432 ) ) - ( $signed( tree_1433 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1437;
always @( posedge clock ) begin
tree_1437 <= ( $signed( tree_1434 ) ) + ( $signed( tree_1435 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1438;
always @( posedge clock ) begin
tree_1438 <=  - ( $signed( tree_1022 ) ) + ( $signed( tree_1024 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1439;
always @( posedge clock ) begin
tree_1439 <= ( $signed( tree_1214 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1440;
always @( posedge clock ) begin
tree_1440 <= ( $signed( tree_1436 ) ) + ( $signed( tree_1437 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1441;
always @( posedge clock ) begin
tree_1441 <= ( $signed( tree_1438 ) ) - ( $signed( tree_1439 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1442;
always @( posedge clock ) begin
tree_1442 <= ( $signed( tree_1440 ) ) + ( $signed( tree_1441 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1443;
always @( posedge clock ) begin
tree_1443 <= ( $signed( in[104] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1444;
always @( posedge clock ) begin
tree_1444 <= ( $signed( tree_1443 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1445;
always @( posedge clock ) begin
tree_1445 <= ( $signed( tree_1444 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1446;
always @( posedge clock ) begin
tree_1446 <= ( $signed( tree_1445 ) ) + ( $signed( tree_1028 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1447;
always @( posedge clock ) begin
tree_1447 <= ( $signed( in[6] ) ) - ( $signed( in[64] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1448;
always @( posedge clock ) begin
tree_1448 <= ( $signed( in[83] ) ) + ( $signed( in[99] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1449;
always @( posedge clock ) begin
tree_1449 <= ( $signed( in[156] ) ) - ( $signed( in[160] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1450;
always @( posedge clock ) begin
tree_1450 <= ( $signed( in[191] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1451;
always @( posedge clock ) begin
tree_1451 <= ( $signed( tree_1447 ) ) - ( $signed( tree_1448 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1452;
always @( posedge clock ) begin
tree_1452 <= ( $signed( tree_1449 ) ) - ( $signed( tree_1450 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1453;
always @( posedge clock ) begin
tree_1453 <= ( $signed( tree_75 ) ) + ( $signed( tree_136 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1454;
always @( posedge clock ) begin
tree_1454 <= ( $signed( tree_326 ) ) + ( $signed( tree_491 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1455;
always @( posedge clock ) begin
tree_1455 <= ( $signed( tree_301 ) ) + ( $signed( tree_456 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1456;
always @( posedge clock ) begin
tree_1456 <= ( $signed( tree_536 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1457;
always @( posedge clock ) begin
tree_1457 <= ( $signed( tree_1451 ) ) + ( $signed( tree_1452 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1458;
always @( posedge clock ) begin
tree_1458 <= ( $signed( tree_1453 ) ) + ( $signed( tree_1454 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1459;
always @( posedge clock ) begin
tree_1459 <=  - ( $signed( tree_1455 ) ) + ( $signed( tree_1456 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1460;
always @( posedge clock ) begin
tree_1460 <= ( $signed( tree_420 ) ) + ( $signed( tree_541 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1461;
always @( posedge clock ) begin
tree_1461 <= ( $signed( tree_543 ) ) + ( $signed( tree_760 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1462;
always @( posedge clock ) begin
tree_1462 <= ( $signed( tree_1457 ) ) - ( $signed( tree_1458 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1463;
always @( posedge clock ) begin
tree_1463 <= ( $signed( tree_1459 ) ) - ( $signed( tree_1460 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1464;
always @( posedge clock ) begin
tree_1464 <= ( $signed( tree_1461 ) ) - ( $signed( tree_1108 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1465;
always @( posedge clock ) begin
tree_1465 <= ( $signed( tree_704 ) ) - ( $signed( tree_836 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1466;
always @( posedge clock ) begin
tree_1466 <= ( $signed( tree_516 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1467;
always @( posedge clock ) begin
tree_1467 <= ( $signed( tree_1462 ) ) + ( $signed( tree_1463 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1468;
always @( posedge clock ) begin
tree_1468 <= ( $signed( tree_1464 ) ) + ( $signed( tree_1465 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1469;
always @( posedge clock ) begin
tree_1469 <= ( $signed( tree_1466 ) ) + ( $signed( tree_1036 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1470;
always @( posedge clock ) begin
tree_1470 <= ( $signed( tree_1467 ) ) + ( $signed( tree_1468 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1471;
always @( posedge clock ) begin
tree_1471 <= ( $signed( tree_1469 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1472;
always @( posedge clock ) begin
tree_1472 <= ( $signed( tree_1470 ) ) - ( $signed( tree_1471 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1473;
always @( posedge clock ) begin
tree_1473 <= ( $signed( in[26] ) ) + ( $signed( in[64] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1474;
always @( posedge clock ) begin
tree_1474 <= ( $signed( in[70] ) ) - ( $signed( in[139] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1475;
always @( posedge clock ) begin
tree_1475 <=  - ( $signed( in[150] ) ) + ( $signed( in[182] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1476;
always @( posedge clock ) begin
tree_1476 <= ( $signed( in[189] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1477;
always @( posedge clock ) begin
tree_1477 <=  - ( $signed( tree_1473 ) ) + ( $signed( tree_1474 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1478;
always @( posedge clock ) begin
tree_1478 <= ( $signed( tree_1475 ) ) + ( $signed( tree_1476 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1479;
always @( posedge clock ) begin
tree_1479 <= ( $signed( tree_30 ) ) + ( $signed( tree_199 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1480;
always @( posedge clock ) begin
tree_1480 <= ( $signed( tree_276 ) ) + ( $signed( tree_138 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1481;
always @( posedge clock ) begin
tree_1481 <=  - ( $signed( tree_323 ) ) + ( $signed( tree_272 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1482;
always @( posedge clock ) begin
tree_1482 <= ( $signed( tree_563 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1483;
always @( posedge clock ) begin
tree_1483 <= ( $signed( tree_1477 ) ) + ( $signed( tree_1478 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1484;
always @( posedge clock ) begin
tree_1484 <=  - ( $signed( tree_1479 ) ) + ( $signed( tree_1480 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1485;
always @( posedge clock ) begin
tree_1485 <= ( $signed( tree_1481 ) ) + ( $signed( tree_1482 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1486;
always @( posedge clock ) begin
tree_1486 <= ( $signed( tree_274 ) ) - ( $signed( tree_724 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1487;
always @( posedge clock ) begin
tree_1487 <= ( $signed( tree_674 ) ) + ( $signed( tree_829 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1488;
always @( posedge clock ) begin
tree_1488 <= ( $signed( tree_822 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1489;
always @( posedge clock ) begin
tree_1489 <= ( $signed( tree_1483 ) ) + ( $signed( tree_1484 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1490;
always @( posedge clock ) begin
tree_1490 <= ( $signed( tree_1485 ) ) + ( $signed( tree_1486 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1491;
always @( posedge clock ) begin
tree_1491 <= ( $signed( tree_1487 ) ) + ( $signed( tree_1488 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1492;
always @( posedge clock ) begin
tree_1492 <= ( $signed( tree_1093 ) ) - ( $signed( tree_1013 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1493;
always @( posedge clock ) begin
tree_1493 <= ( $signed( tree_1041 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1494;
always @( posedge clock ) begin
tree_1494 <= ( $signed( tree_1489 ) ) + ( $signed( tree_1490 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1495;
always @( posedge clock ) begin
tree_1495 <=  - ( $signed( tree_1491 ) ) + ( $signed( tree_1492 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1496;
always @( posedge clock ) begin
tree_1496 <= ( $signed( tree_1493 ) ) + ( $signed( tree_1276 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1497;
always @( posedge clock ) begin
tree_1497 <= ( $signed( tree_1494 ) ) + ( $signed( tree_1495 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1498;
always @( posedge clock ) begin
tree_1498 <= ( $signed( tree_1496 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1499;
always @( posedge clock ) begin
tree_1499 <= ( $signed( tree_1497 ) ) - ( $signed( tree_1498 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1500;
always @( posedge clock ) begin
tree_1500 <= ( $signed( in[61] ) ) - ( $signed( in[85] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1501;
always @( posedge clock ) begin
tree_1501 <= ( $signed( in[93] ) ) + ( $signed( in[108] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1502;
always @( posedge clock ) begin
tree_1502 <= ( $signed( in[155] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1503;
always @( posedge clock ) begin
tree_1503 <= ( $signed( tree_1500 ) ) + ( $signed( tree_1501 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1504;
always @( posedge clock ) begin
tree_1504 <= ( $signed( tree_1502 ) ) + ( $signed( tree_75 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1505;
always @( posedge clock ) begin
tree_1505 <=  - ( $signed( tree_146 ) ) + ( $signed( tree_210 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1506;
always @( posedge clock ) begin
tree_1506 <= ( $signed( tree_20 ) ) - ( $signed( tree_398 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1507;
always @( posedge clock ) begin
tree_1507 <= ( $signed( tree_568 ) ) + ( $signed( tree_455 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1508;
always @( posedge clock ) begin
tree_1508 <= ( $signed( tree_8 ) ) + ( $signed( tree_461 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1509;
always @( posedge clock ) begin
tree_1509 <= ( $signed( tree_571 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1510;
always @( posedge clock ) begin
tree_1510 <= ( $signed( tree_1503 ) ) + ( $signed( tree_1504 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1511;
always @( posedge clock ) begin
tree_1511 <= ( $signed( tree_1505 ) ) + ( $signed( tree_1506 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1512;
always @( posedge clock ) begin
tree_1512 <= ( $signed( tree_1507 ) ) + ( $signed( tree_1508 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1513;
always @( posedge clock ) begin
tree_1513 <= ( $signed( tree_1509 ) ) + ( $signed( tree_361 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1514;
always @( posedge clock ) begin
tree_1514 <= ( $signed( tree_212 ) ) - ( $signed( tree_443 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1515;
always @( posedge clock ) begin
tree_1515 <= ( $signed( tree_497 ) ) + ( $signed( tree_570 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1516;
always @( posedge clock ) begin
tree_1516 <= ( $signed( tree_572 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1517;
always @( posedge clock ) begin
tree_1517 <= ( $signed( tree_1510 ) ) + ( $signed( tree_1511 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1518;
always @( posedge clock ) begin
tree_1518 <= ( $signed( tree_1512 ) ) + ( $signed( tree_1513 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1519;
always @( posedge clock ) begin
tree_1519 <= ( $signed( tree_1514 ) ) - ( $signed( tree_1515 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1520;
always @( posedge clock ) begin
tree_1520 <= ( $signed( tree_1516 ) ) + ( $signed( tree_939 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1521;
always @( posedge clock ) begin
tree_1521 <= ( $signed( tree_989 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1522;
always @( posedge clock ) begin
tree_1522 <= ( $signed( tree_1517 ) ) - ( $signed( tree_1518 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1523;
always @( posedge clock ) begin
tree_1523 <= ( $signed( tree_1519 ) ) + ( $signed( tree_1520 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1524;
always @( posedge clock ) begin
tree_1524 <= ( $signed( tree_1521 ) ) + ( $signed( tree_1189 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1525;
always @( posedge clock ) begin
tree_1525 <= ( $signed( tree_1522 ) ) + ( $signed( tree_1523 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1526;
always @( posedge clock ) begin
tree_1526 <= ( $signed( tree_1524 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1527;
always @( posedge clock ) begin
tree_1527 <= ( $signed( tree_1525 ) ) + ( $signed( tree_1526 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1528;
always @( posedge clock ) begin
tree_1528 <= ( $signed( tree_80 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1529;
always @( posedge clock ) begin
tree_1529 <= ( $signed( tree_1528 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1530;
always @( posedge clock ) begin
tree_1530 <= ( $signed( tree_1529 ) ) - ( $signed( tree_1141 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1531;
always @( posedge clock ) begin
tree_1531 <= ( $signed( in[29] ) ) + ( $signed( in[102] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1532;
always @( posedge clock ) begin
tree_1532 <= ( $signed( in[175] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1533;
always @( posedge clock ) begin
tree_1533 <=  - ( $signed( tree_1531 ) ) + ( $signed( tree_1532 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1534;
always @( posedge clock ) begin
tree_1534 <=  - ( $signed( tree_9 ) ) + ( $signed( tree_17 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1535;
always @( posedge clock ) begin
tree_1535 <= ( $signed( tree_142 ) ) + ( $signed( tree_134 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1536;
always @( posedge clock ) begin
tree_1536 <= ( $signed( tree_296 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1537;
always @( posedge clock ) begin
tree_1537 <= ( $signed( tree_1533 ) ) + ( $signed( tree_1534 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1538;
always @( posedge clock ) begin
tree_1538 <= ( $signed( tree_1535 ) ) + ( $signed( tree_1536 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1539;
always @( posedge clock ) begin
tree_1539 <=  - ( $signed( tree_774 ) ) + ( $signed( tree_723 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1540;
always @( posedge clock ) begin
tree_1540 <= ( $signed( tree_558 ) ) - ( $signed( tree_583 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1541;
always @( posedge clock ) begin
tree_1541 <= ( $signed( tree_806 ) ) + ( $signed( tree_837 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1542;
always @( posedge clock ) begin
tree_1542 <= ( $signed( tree_1047 ) ) - ( $signed( tree_575 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1543;
always @( posedge clock ) begin
tree_1543 <= ( $signed( tree_460 ) ) + ( $signed( tree_587 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1544;
always @( posedge clock ) begin
tree_1544 <= ( $signed( tree_1537 ) ) + ( $signed( tree_1538 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1545;
always @( posedge clock ) begin
tree_1545 <= ( $signed( tree_1539 ) ) + ( $signed( tree_1540 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1546;
always @( posedge clock ) begin
tree_1546 <=  - ( $signed( tree_1541 ) ) + ( $signed( tree_1542 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1547;
always @( posedge clock ) begin
tree_1547 <= ( $signed( tree_1543 ) ) + ( $signed( tree_1100 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1548;
always @( posedge clock ) begin
tree_1548 <=  - ( $signed( tree_581 ) ) + ( $signed( tree_848 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1549;
always @( posedge clock ) begin
tree_1549 <= ( $signed( tree_384 ) ) + ( $signed( tree_1049 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1550;
always @( posedge clock ) begin
tree_1550 <= ( $signed( tree_970 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1551;
always @( posedge clock ) begin
tree_1551 <= ( $signed( tree_1544 ) ) + ( $signed( tree_1545 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1552;
always @( posedge clock ) begin
tree_1552 <= ( $signed( tree_1546 ) ) + ( $signed( tree_1547 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1553;
always @( posedge clock ) begin
tree_1553 <= ( $signed( tree_1548 ) ) - ( $signed( tree_1549 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1554;
always @( posedge clock ) begin
tree_1554 <= ( $signed( tree_1550 ) ) + ( $signed( tree_964 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1555;
always @( posedge clock ) begin
tree_1555 <= ( $signed( tree_1551 ) ) + ( $signed( tree_1552 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1556;
always @( posedge clock ) begin
tree_1556 <= ( $signed( tree_1553 ) ) - ( $signed( tree_1554 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1557;
always @( posedge clock ) begin
tree_1557 <= ( $signed( tree_1555 ) ) + ( $signed( tree_1556 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1558;
always @( posedge clock ) begin
tree_1558 <= ( $signed( in[109] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1559;
always @( posedge clock ) begin
tree_1559 <= ( $signed( tree_1558 ) ) - ( $signed( tree_199 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1560;
always @( posedge clock ) begin
tree_1560 <= ( $signed( tree_188 ) ) + ( $signed( tree_189 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1561;
always @( posedge clock ) begin
tree_1561 <= ( $signed( tree_126 ) ) - ( $signed( tree_518 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1562;
always @( posedge clock ) begin
tree_1562 <=  - ( $signed( tree_201 ) ) + ( $signed( tree_498 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1563;
always @( posedge clock ) begin
tree_1563 <= ( $signed( tree_588 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1564;
always @( posedge clock ) begin
tree_1564 <= ( $signed( tree_1559 ) ) - ( $signed( tree_1560 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1565;
always @( posedge clock ) begin
tree_1565 <= ( $signed( tree_1561 ) ) + ( $signed( tree_1562 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1566;
always @( posedge clock ) begin
tree_1566 <= ( $signed( tree_1563 ) ) + ( $signed( tree_776 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1567;
always @( posedge clock ) begin
tree_1567 <= ( $signed( tree_111 ) ) + ( $signed( tree_393 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1568;
always @( posedge clock ) begin
tree_1568 <= ( $signed( tree_646 ) ) - ( $signed( tree_547 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1569;
always @( posedge clock ) begin
tree_1569 <= ( $signed( tree_1564 ) ) + ( $signed( tree_1565 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1570;
always @( posedge clock ) begin
tree_1570 <=  - ( $signed( tree_1566 ) ) + ( $signed( tree_1567 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1571;
always @( posedge clock ) begin
tree_1571 <= ( $signed( tree_1568 ) ) - ( $signed( tree_832 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1572;
always @( posedge clock ) begin
tree_1572 <=  - ( $signed( tree_1052 ) ) + ( $signed( tree_995 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1573;
always @( posedge clock ) begin
tree_1573 <= ( $signed( tree_748 ) ) - ( $signed( tree_1017 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1574;
always @( posedge clock ) begin
tree_1574 <= ( $signed( tree_1178 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1575;
always @( posedge clock ) begin
tree_1575 <= ( $signed( tree_1569 ) ) + ( $signed( tree_1570 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1576;
always @( posedge clock ) begin
tree_1576 <= ( $signed( tree_1571 ) ) + ( $signed( tree_1572 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1577;
always @( posedge clock ) begin
tree_1577 <= ( $signed( tree_1573 ) ) - ( $signed( tree_1574 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1578;
always @( posedge clock ) begin
tree_1578 <= ( $signed( tree_1022 ) ) + ( $signed( tree_1054 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1579;
always @( posedge clock ) begin
tree_1579 <= ( $signed( tree_1575 ) ) + ( $signed( tree_1576 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1580;
always @( posedge clock ) begin
tree_1580 <= ( $signed( tree_1577 ) ) - ( $signed( tree_1578 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1581;
always @( posedge clock ) begin
tree_1581 <= ( $signed( tree_1058 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1582;
always @( posedge clock ) begin
tree_1582 <= ( $signed( tree_1579 ) ) + ( $signed( tree_1580 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1583;
always @( posedge clock ) begin
tree_1583 <= ( $signed( tree_1581 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1584;
always @( posedge clock ) begin
tree_1584 <= ( $signed( tree_1582 ) ) + ( $signed( tree_1583 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1585;
always @( posedge clock ) begin
tree_1585 <= ( $signed( tree_121 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1586;
always @( posedge clock ) begin
tree_1586 <= ( $signed( tree_1585 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1587;
always @( posedge clock ) begin
tree_1587 <= ( $signed( tree_1586 ) ) - ( $signed( tree_1119 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1588;
always @( posedge clock ) begin
tree_1588 <= ( $signed( in[6] ) ) + ( $signed( in[102] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1589;
always @( posedge clock ) begin
tree_1589 <=  - ( $signed( in[155] ) ) + ( $signed( in[167] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1590;
always @( posedge clock ) begin
tree_1590 <=  - ( $signed( tree_1588 ) ) + ( $signed( tree_1589 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1591;
always @( posedge clock ) begin
tree_1591 <= ( $signed( tree_99 ) ) + ( $signed( tree_61 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1592;
always @( posedge clock ) begin
tree_1592 <= ( $signed( tree_319 ) ) + ( $signed( tree_376 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1593;
always @( posedge clock ) begin
tree_1593 <= ( $signed( tree_601 ) ) - ( $signed( tree_374 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1594;
always @( posedge clock ) begin
tree_1594 <= ( $signed( tree_333 ) ) + ( $signed( tree_469 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1595;
always @( posedge clock ) begin
tree_1595 <= ( $signed( tree_251 ) ) - ( $signed( tree_602 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1596;
always @( posedge clock ) begin
tree_1596 <= ( $signed( tree_1590 ) ) + ( $signed( tree_1591 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1597;
always @( posedge clock ) begin
tree_1597 <= ( $signed( tree_1592 ) ) + ( $signed( tree_1593 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1598;
always @( posedge clock ) begin
tree_1598 <= ( $signed( tree_1594 ) ) + ( $signed( tree_1595 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1599;
always @( posedge clock ) begin
tree_1599 <= ( $signed( tree_692 ) ) - ( $signed( tree_463 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1600;
always @( posedge clock ) begin
tree_1600 <= ( $signed( tree_267 ) ) - ( $signed( tree_128 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1601;
always @( posedge clock ) begin
tree_1601 <= ( $signed( tree_429 ) ) + ( $signed( tree_347 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1602;
always @( posedge clock ) begin
tree_1602 <=  - ( $signed( tree_570 ) ) + ( $signed( tree_1014 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1603;
always @( posedge clock ) begin
tree_1603 <= ( $signed( tree_579 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1604;
always @( posedge clock ) begin
tree_1604 <= ( $signed( tree_1596 ) ) + ( $signed( tree_1597 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1605;
always @( posedge clock ) begin
tree_1605 <= ( $signed( tree_1598 ) ) + ( $signed( tree_1599 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1606;
always @( posedge clock ) begin
tree_1606 <= ( $signed( tree_1600 ) ) + ( $signed( tree_1601 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1607;
always @( posedge clock ) begin
tree_1607 <= ( $signed( tree_1602 ) ) + ( $signed( tree_1603 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1608;
always @( posedge clock ) begin
tree_1608 <= ( $signed( tree_874 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1609;
always @( posedge clock ) begin
tree_1609 <= ( $signed( tree_1604 ) ) + ( $signed( tree_1605 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1610;
always @( posedge clock ) begin
tree_1610 <= ( $signed( tree_1606 ) ) + ( $signed( tree_1607 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1611;
always @( posedge clock ) begin
tree_1611 <=  - ( $signed( tree_1608 ) ) + ( $signed( tree_1174 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1612;
always @( posedge clock ) begin
tree_1612 <= ( $signed( tree_1609 ) ) + ( $signed( tree_1610 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1613;
always @( posedge clock ) begin
tree_1613 <= ( $signed( tree_1611 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1614;
always @( posedge clock ) begin
tree_1614 <= ( $signed( tree_1612 ) ) + ( $signed( tree_1613 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1615;
always @( posedge clock ) begin
tree_1615 <= ( $signed( tree_254 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1616;
always @( posedge clock ) begin
tree_1616 <= ( $signed( tree_1615 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1617;
always @( posedge clock ) begin
tree_1617 <= ( $signed( tree_1616 ) ) + ( $signed( tree_1060 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1618;
always @( posedge clock ) begin
tree_1618 <= ( $signed( in[2] ) ) + ( $signed( in[40] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1619;
always @( posedge clock ) begin
tree_1619 <= ( $signed( in[110] ) ) + ( $signed( in[132] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1620;
always @( posedge clock ) begin
tree_1620 <= ( $signed( in[133] ) ) + ( $signed( in[154] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1621;
always @( posedge clock ) begin
tree_1621 <= ( $signed( in[156] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1622;
always @( posedge clock ) begin
tree_1622 <= ( $signed( tree_1618 ) ) + ( $signed( tree_1619 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1623;
always @( posedge clock ) begin
tree_1623 <= ( $signed( tree_1620 ) ) + ( $signed( tree_1621 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1624;
always @( posedge clock ) begin
tree_1624 <= ( $signed( tree_13 ) ) + ( $signed( tree_265 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1625;
always @( posedge clock ) begin
tree_1625 <= ( $signed( tree_408 ) ) + ( $signed( tree_601 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1626;
always @( posedge clock ) begin
tree_1626 <=  - ( $signed( tree_134 ) ) + ( $signed( tree_194 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1627;
always @( posedge clock ) begin
tree_1627 <= ( $signed( tree_617 ) ) + ( $signed( tree_618 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1628;
always @( posedge clock ) begin
tree_1628 <= ( $signed( tree_1622 ) ) + ( $signed( tree_1623 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1629;
always @( posedge clock ) begin
tree_1629 <= ( $signed( tree_1624 ) ) + ( $signed( tree_1625 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1630;
always @( posedge clock ) begin
tree_1630 <= ( $signed( tree_1626 ) ) + ( $signed( tree_1627 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1631;
always @( posedge clock ) begin
tree_1631 <= ( $signed( tree_701 ) ) + ( $signed( tree_952 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1632;
always @( posedge clock ) begin
tree_1632 <=  - ( $signed( tree_665 ) ) + ( $signed( tree_468 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1633;
always @( posedge clock ) begin
tree_1633 <=  - ( $signed( tree_583 ) ) + ( $signed( tree_431 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1634;
always @( posedge clock ) begin
tree_1634 <=  - ( $signed( tree_1628 ) ) + ( $signed( tree_1629 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1635;
always @( posedge clock ) begin
tree_1635 <= ( $signed( tree_1630 ) ) + ( $signed( tree_1631 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1636;
always @( posedge clock ) begin
tree_1636 <= ( $signed( tree_1632 ) ) + ( $signed( tree_1633 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1637;
always @( posedge clock ) begin
tree_1637 <= ( $signed( tree_851 ) ) - ( $signed( tree_574 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1638;
always @( posedge clock ) begin
tree_1638 <= ( $signed( tree_903 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1639;
always @( posedge clock ) begin
tree_1639 <= ( $signed( tree_1634 ) ) + ( $signed( tree_1635 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1640;
always @( posedge clock ) begin
tree_1640 <= ( $signed( tree_1636 ) ) + ( $signed( tree_1637 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1641;
always @( posedge clock ) begin
tree_1641 <= ( $signed( tree_1638 ) ) - ( $signed( tree_993 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1642;
always @( posedge clock ) begin
tree_1642 <= ( $signed( tree_1062 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1643;
always @( posedge clock ) begin
tree_1643 <= ( $signed( tree_1639 ) ) + ( $signed( tree_1640 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1644;
always @( posedge clock ) begin
tree_1644 <= ( $signed( tree_1641 ) ) - ( $signed( tree_1642 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1645;
always @( posedge clock ) begin
tree_1645 <= ( $signed( tree_1643 ) ) + ( $signed( tree_1644 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1646;
always @( posedge clock ) begin
tree_1646 <= ( $signed( in[19] ) ) + ( $signed( in[21] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1647;
always @( posedge clock ) begin
tree_1647 <= ( $signed( in[108] ) ) + ( $signed( in[130] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1648;
always @( posedge clock ) begin
tree_1648 <= ( $signed( in[178] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1649;
always @( posedge clock ) begin
tree_1649 <= ( $signed( tree_1646 ) ) + ( $signed( tree_1647 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1650;
always @( posedge clock ) begin
tree_1650 <=  - ( $signed( tree_1648 ) ) + ( $signed( tree_162 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1651;
always @( posedge clock ) begin
tree_1651 <= ( $signed( tree_202 ) ) + ( $signed( tree_60 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1652;
always @( posedge clock ) begin
tree_1652 <= ( $signed( tree_225 ) ) - ( $signed( tree_264 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1653;
always @( posedge clock ) begin
tree_1653 <= ( $signed( tree_341 ) ) + ( $signed( tree_198 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1654;
always @( posedge clock ) begin
tree_1654 <= ( $signed( tree_490 ) ) + ( $signed( tree_190 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1655;
always @( posedge clock ) begin
tree_1655 <= ( $signed( tree_230 ) ) + ( $signed( tree_233 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1656;
always @( posedge clock ) begin
tree_1656 <= ( $signed( tree_108 ) ) + ( $signed( tree_521 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1657;
always @( posedge clock ) begin
tree_1657 <= ( $signed( tree_1649 ) ) + ( $signed( tree_1650 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1658;
always @( posedge clock ) begin
tree_1658 <=  - ( $signed( tree_1651 ) ) + ( $signed( tree_1652 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1659;
always @( posedge clock ) begin
tree_1659 <= ( $signed( tree_1653 ) ) + ( $signed( tree_1654 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1660;
always @( posedge clock ) begin
tree_1660 <= ( $signed( tree_1655 ) ) + ( $signed( tree_1656 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1661;
always @( posedge clock ) begin
tree_1661 <=  - ( $signed( tree_808 ) ) + ( $signed( tree_375 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1662;
always @( posedge clock ) begin
tree_1662 <= ( $signed( tree_178 ) ) - ( $signed( tree_927 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1663;
always @( posedge clock ) begin
tree_1663 <= ( $signed( tree_870 ) ) + ( $signed( tree_943 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1664;
always @( posedge clock ) begin
tree_1664 <= ( $signed( tree_1657 ) ) + ( $signed( tree_1658 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1665;
always @( posedge clock ) begin
tree_1665 <= ( $signed( tree_1659 ) ) + ( $signed( tree_1660 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1666;
always @( posedge clock ) begin
tree_1666 <= ( $signed( tree_1661 ) ) + ( $signed( tree_1662 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1667;
always @( posedge clock ) begin
tree_1667 <=  - ( $signed( tree_1663 ) ) + ( $signed( tree_524 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1668;
always @( posedge clock ) begin
tree_1668 <= ( $signed( tree_1165 ) ) + ( $signed( tree_399 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1669;
always @( posedge clock ) begin
tree_1669 <= ( $signed( tree_1664 ) ) + ( $signed( tree_1665 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1670;
always @( posedge clock ) begin
tree_1670 <= ( $signed( tree_1666 ) ) + ( $signed( tree_1667 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1671;
always @( posedge clock ) begin
tree_1671 <= ( $signed( tree_1668 ) ) - ( $signed( tree_1223 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1672;
always @( posedge clock ) begin
tree_1672 <= ( $signed( tree_1669 ) ) + ( $signed( tree_1670 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1673;
always @( posedge clock ) begin
tree_1673 <= ( $signed( tree_1671 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1674;
always @( posedge clock ) begin
tree_1674 <= ( $signed( tree_1672 ) ) + ( $signed( tree_1673 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1675;
always @( posedge clock ) begin
tree_1675 <= ( $signed( in[50] ) ) - ( $signed( in[167] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1676;
always @( posedge clock ) begin
tree_1676 <= ( $signed( tree_1675 ) ) - ( $signed( tree_76 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1677;
always @( posedge clock ) begin
tree_1677 <= ( $signed( tree_64 ) ) + ( $signed( tree_307 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1678;
always @( posedge clock ) begin
tree_1678 <= ( $signed( tree_454 ) ) - ( $signed( tree_588 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1679;
always @( posedge clock ) begin
tree_1679 <= ( $signed( tree_1676 ) ) - ( $signed( tree_1677 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1680;
always @( posedge clock ) begin
tree_1680 <= ( $signed( tree_1678 ) ) - ( $signed( tree_106 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1681;
always @( posedge clock ) begin
tree_1681 <= ( $signed( tree_91 ) ) + ( $signed( tree_854 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1682;
always @( posedge clock ) begin
tree_1682 <=  - ( $signed( tree_423 ) ) + ( $signed( tree_459 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1683;
always @( posedge clock ) begin
tree_1683 <= ( $signed( tree_764 ) ) - ( $signed( tree_661 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1684;
always @( posedge clock ) begin
tree_1684 <= ( $signed( tree_875 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1685;
always @( posedge clock ) begin
tree_1685 <= ( $signed( tree_1679 ) ) + ( $signed( tree_1680 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1686;
always @( posedge clock ) begin
tree_1686 <=  - ( $signed( tree_1681 ) ) + ( $signed( tree_1682 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1687;
always @( posedge clock ) begin
tree_1687 <= ( $signed( tree_1683 ) ) + ( $signed( tree_1684 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1688;
always @( posedge clock ) begin
tree_1688 <= ( $signed( tree_1202 ) ) - ( $signed( tree_608 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1689;
always @( posedge clock ) begin
tree_1689 <= ( $signed( tree_1103 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1690;
always @( posedge clock ) begin
tree_1690 <= ( $signed( tree_1685 ) ) + ( $signed( tree_1686 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1691;
always @( posedge clock ) begin
tree_1691 <= ( $signed( tree_1687 ) ) + ( $signed( tree_1688 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1692;
always @( posedge clock ) begin
tree_1692 <= ( $signed( tree_1689 ) ) + ( $signed( tree_1024 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1693;
always @( posedge clock ) begin
tree_1693 <= ( $signed( tree_1690 ) ) + ( $signed( tree_1691 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1694;
always @( posedge clock ) begin
tree_1694 <= ( $signed( tree_1692 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1695;
always @( posedge clock ) begin
tree_1695 <= ( $signed( tree_1693 ) ) + ( $signed( tree_1694 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1696;
always @( posedge clock ) begin
tree_1696 <= ( $signed( in[10] ) ) + ( $signed( in[59] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1697;
always @( posedge clock ) begin
tree_1697 <= ( $signed( in[88] ) ) + ( $signed( in[106] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1698;
always @( posedge clock ) begin
tree_1698 <= ( $signed( in[114] ) ) + ( $signed( in[115] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1699;
always @( posedge clock ) begin
tree_1699 <=  - ( $signed( in[123] ) ) + ( $signed( in[150] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1700;
always @( posedge clock ) begin
tree_1700 <= ( $signed( tree_1696 ) ) - ( $signed( tree_1697 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1701;
always @( posedge clock ) begin
tree_1701 <=  - ( $signed( tree_1698 ) ) + ( $signed( tree_1699 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1702;
always @( posedge clock ) begin
tree_1702 <= ( $signed( tree_27 ) ) + ( $signed( tree_331 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1703;
always @( posedge clock ) begin
tree_1703 <= ( $signed( tree_149 ) ) + ( $signed( tree_301 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1704;
always @( posedge clock ) begin
tree_1704 <= ( $signed( tree_329 ) ) + ( $signed( tree_467 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1705;
always @( posedge clock ) begin
tree_1705 <= ( $signed( tree_502 ) ) - ( $signed( tree_584 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1706;
always @( posedge clock ) begin
tree_1706 <= ( $signed( tree_571 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1707;
always @( posedge clock ) begin
tree_1707 <= ( $signed( tree_1700 ) ) + ( $signed( tree_1701 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1708;
always @( posedge clock ) begin
tree_1708 <= ( $signed( tree_1702 ) ) + ( $signed( tree_1703 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1709;
always @( posedge clock ) begin
tree_1709 <=  - ( $signed( tree_1704 ) ) + ( $signed( tree_1705 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1710;
always @( posedge clock ) begin
tree_1710 <= ( $signed( tree_1706 ) ) + ( $signed( tree_363 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1711;
always @( posedge clock ) begin
tree_1711 <=  - ( $signed( tree_647 ) ) + ( $signed( tree_594 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1712;
always @( posedge clock ) begin
tree_1712 <= ( $signed( tree_746 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1713;
always @( posedge clock ) begin
tree_1713 <= ( $signed( tree_1707 ) ) - ( $signed( tree_1708 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1714;
always @( posedge clock ) begin
tree_1714 <= ( $signed( tree_1709 ) ) - ( $signed( tree_1710 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1715;
always @( posedge clock ) begin
tree_1715 <= ( $signed( tree_1711 ) ) + ( $signed( tree_1712 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1716;
always @( posedge clock ) begin
tree_1716 <= ( $signed( tree_1006 ) ) + ( $signed( tree_505 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1717;
always @( posedge clock ) begin
tree_1717 <= ( $signed( tree_1713 ) ) + ( $signed( tree_1714 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1718;
always @( posedge clock ) begin
tree_1718 <= ( $signed( tree_1715 ) ) + ( $signed( tree_1716 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1719;
always @( posedge clock ) begin
tree_1719 <= ( $signed( tree_1530 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1720;
always @( posedge clock ) begin
tree_1720 <= ( $signed( tree_1717 ) ) + ( $signed( tree_1718 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1721;
always @( posedge clock ) begin
tree_1721 <= ( $signed( tree_1719 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1722;
always @( posedge clock ) begin
tree_1722 <= ( $signed( tree_1720 ) ) + ( $signed( tree_1721 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1723;
always @( posedge clock ) begin
tree_1723 <= ( $signed( in[24] ) ) - ( $signed( in[33] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1724;
always @( posedge clock ) begin
tree_1724 <= ( $signed( tree_1723 ) ) + ( $signed( tree_18 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1725;
always @( posedge clock ) begin
tree_1725 <= ( $signed( tree_118 ) ) + ( $signed( tree_2 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1726;
always @( posedge clock ) begin
tree_1726 <= ( $signed( tree_163 ) ) + ( $signed( tree_601 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1727;
always @( posedge clock ) begin
tree_1727 <= ( $signed( tree_221 ) ) + ( $signed( tree_626 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1728;
always @( posedge clock ) begin
tree_1728 <= ( $signed( tree_627 ) ) - ( $signed( tree_421 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1729;
always @( posedge clock ) begin
tree_1729 <= ( $signed( tree_1724 ) ) + ( $signed( tree_1725 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1730;
always @( posedge clock ) begin
tree_1730 <= ( $signed( tree_1726 ) ) + ( $signed( tree_1727 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1731;
always @( posedge clock ) begin
tree_1731 <= ( $signed( tree_1728 ) ) + ( $signed( tree_340 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1732;
always @( posedge clock ) begin
tree_1732 <= ( $signed( tree_159 ) ) - ( $signed( tree_155 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1733;
always @( posedge clock ) begin
tree_1733 <=  - ( $signed( tree_629 ) ) + ( $signed( tree_1047 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1734;
always @( posedge clock ) begin
tree_1734 <= ( $signed( tree_612 ) ) + ( $signed( tree_1019 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1735;
always @( posedge clock ) begin
tree_1735 <= ( $signed( tree_1729 ) ) - ( $signed( tree_1730 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1736;
always @( posedge clock ) begin
tree_1736 <= ( $signed( tree_1731 ) ) + ( $signed( tree_1732 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1737;
always @( posedge clock ) begin
tree_1737 <= ( $signed( tree_1733 ) ) + ( $signed( tree_1734 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1738;
always @( posedge clock ) begin
tree_1738 <= ( $signed( tree_1260 ) ) - ( $signed( tree_535 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1739;
always @( posedge clock ) begin
tree_1739 <= ( $signed( tree_987 ) ) + ( $signed( tree_1002 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1740;
always @( posedge clock ) begin
tree_1740 <= ( $signed( tree_766 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1741;
always @( posedge clock ) begin
tree_1741 <= ( $signed( tree_1735 ) ) + ( $signed( tree_1736 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1742;
always @( posedge clock ) begin
tree_1742 <= ( $signed( tree_1737 ) ) + ( $signed( tree_1738 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1743;
always @( posedge clock ) begin
tree_1743 <= ( $signed( tree_1739 ) ) + ( $signed( tree_1740 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1744;
always @( posedge clock ) begin
tree_1744 <= ( $signed( tree_1036 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1745;
always @( posedge clock ) begin
tree_1745 <= ( $signed( tree_1741 ) ) + ( $signed( tree_1742 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1746;
always @( posedge clock ) begin
tree_1746 <= ( $signed( tree_1743 ) ) + ( $signed( tree_1744 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1747;
always @( posedge clock ) begin
tree_1747 <= ( $signed( tree_1745 ) ) + ( $signed( tree_1746 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1748;
always @( posedge clock ) begin
tree_1748 <= ( $signed( in[12] ) ) - ( $signed( in[17] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1749;
always @( posedge clock ) begin
tree_1749 <= ( $signed( in[51] ) ) - ( $signed( in[78] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1750;
always @( posedge clock ) begin
tree_1750 <= ( $signed( in[86] ) ) + ( $signed( in[120] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1751;
always @( posedge clock ) begin
tree_1751 <= ( $signed( in[165] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1752;
always @( posedge clock ) begin
tree_1752 <= ( $signed( tree_1748 ) ) + ( $signed( tree_1749 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1753;
always @( posedge clock ) begin
tree_1753 <= ( $signed( tree_1750 ) ) + ( $signed( tree_1751 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1754;
always @( posedge clock ) begin
tree_1754 <=  - ( $signed( tree_40 ) ) + ( $signed( tree_88 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1755;
always @( posedge clock ) begin
tree_1755 <= ( $signed( tree_93 ) ) - ( $signed( tree_24 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1756;
always @( posedge clock ) begin
tree_1756 <= ( $signed( tree_168 ) ) + ( $signed( tree_416 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1757;
always @( posedge clock ) begin
tree_1757 <= ( $signed( tree_467 ) ) + ( $signed( tree_626 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1758;
always @( posedge clock ) begin
tree_1758 <=  - ( $signed( tree_480 ) ) + ( $signed( tree_602 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1759;
always @( posedge clock ) begin
tree_1759 <= ( $signed( tree_1752 ) ) - ( $signed( tree_1753 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1760;
always @( posedge clock ) begin
tree_1760 <= ( $signed( tree_1754 ) ) + ( $signed( tree_1755 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1761;
always @( posedge clock ) begin
tree_1761 <= ( $signed( tree_1756 ) ) - ( $signed( tree_1757 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1762;
always @( posedge clock ) begin
tree_1762 <= ( $signed( tree_1758 ) ) - ( $signed( tree_565 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1763;
always @( posedge clock ) begin
tree_1763 <= ( $signed( tree_629 ) ) + ( $signed( tree_572 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1764;
always @( posedge clock ) begin
tree_1764 <= ( $signed( tree_1759 ) ) + ( $signed( tree_1760 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1765;
always @( posedge clock ) begin
tree_1765 <= ( $signed( tree_1761 ) ) + ( $signed( tree_1762 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1766;
always @( posedge clock ) begin
tree_1766 <= ( $signed( tree_1763 ) ) + ( $signed( tree_865 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1767;
always @( posedge clock ) begin
tree_1767 <= ( $signed( tree_1098 ) ) + ( $signed( tree_219 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1768;
always @( posedge clock ) begin
tree_1768 <=  - ( $signed( tree_986 ) ) + ( $signed( tree_1177 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1769;
always @( posedge clock ) begin
tree_1769 <= ( $signed( tree_1764 ) ) + ( $signed( tree_1765 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1770;
always @( posedge clock ) begin
tree_1770 <= ( $signed( tree_1766 ) ) + ( $signed( tree_1767 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1771;
always @( posedge clock ) begin
tree_1771 <= ( $signed( tree_1768 ) ) - ( $signed( tree_1266 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1772;
always @( posedge clock ) begin
tree_1772 <= ( $signed( tree_1043 ) ) + ( $signed( tree_1088 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1773;
always @( posedge clock ) begin
tree_1773 <= ( $signed( tree_1769 ) ) + ( $signed( tree_1770 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1774;
always @( posedge clock ) begin
tree_1774 <= ( $signed( tree_1771 ) ) - ( $signed( tree_1772 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1775;
always @( posedge clock ) begin
tree_1775 <= ( $signed( tree_1773 ) ) + ( $signed( tree_1774 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1776;
always @( posedge clock ) begin
tree_1776 <= ( $signed( in[135] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1777;
always @( posedge clock ) begin
tree_1777 <= ( $signed( tree_1776 ) ) + ( $signed( tree_33 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1778;
always @( posedge clock ) begin
tree_1778 <= ( $signed( tree_147 ) ) + ( $signed( tree_202 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1779;
always @( posedge clock ) begin
tree_1779 <=  - ( $signed( tree_189 ) ) + ( $signed( tree_169 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1780;
always @( posedge clock ) begin
tree_1780 <= ( $signed( tree_113 ) ) + ( $signed( tree_333 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1781;
always @( posedge clock ) begin
tree_1781 <=  - ( $signed( tree_627 ) ) + ( $signed( tree_501 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1782;
always @( posedge clock ) begin
tree_1782 <= ( $signed( tree_563 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1783;
always @( posedge clock ) begin
tree_1783 <= ( $signed( tree_1777 ) ) + ( $signed( tree_1778 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1784;
always @( posedge clock ) begin
tree_1784 <= ( $signed( tree_1779 ) ) - ( $signed( tree_1780 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1785;
always @( posedge clock ) begin
tree_1785 <= ( $signed( tree_1781 ) ) - ( $signed( tree_1782 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1786;
always @( posedge clock ) begin
tree_1786 <= ( $signed( tree_259 ) ) + ( $signed( tree_171 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1787;
always @( posedge clock ) begin
tree_1787 <= ( $signed( tree_285 ) ) + ( $signed( tree_500 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1788;
always @( posedge clock ) begin
tree_1788 <= ( $signed( tree_433 ) ) + ( $signed( tree_911 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1789;
always @( posedge clock ) begin
tree_1789 <= ( $signed( tree_616 ) ) + ( $signed( tree_631 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1790;
always @( posedge clock ) begin
tree_1790 <= ( $signed( tree_757 ) ) + ( $signed( tree_936 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1791;
always @( posedge clock ) begin
tree_1791 <= ( $signed( tree_587 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1792;
always @( posedge clock ) begin
tree_1792 <=  - ( $signed( tree_1783 ) ) + ( $signed( tree_1784 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1793;
always @( posedge clock ) begin
tree_1793 <= ( $signed( tree_1785 ) ) - ( $signed( tree_1786 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1794;
always @( posedge clock ) begin
tree_1794 <= ( $signed( tree_1787 ) ) + ( $signed( tree_1788 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1795;
always @( posedge clock ) begin
tree_1795 <= ( $signed( tree_1789 ) ) + ( $signed( tree_1790 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1796;
always @( posedge clock ) begin
tree_1796 <=  - ( $signed( tree_1791 ) ) + ( $signed( tree_611 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1797;
always @( posedge clock ) begin
tree_1797 <= ( $signed( tree_1264 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1798;
always @( posedge clock ) begin
tree_1798 <= ( $signed( tree_1792 ) ) + ( $signed( tree_1793 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1799;
always @( posedge clock ) begin
tree_1799 <= ( $signed( tree_1794 ) ) + ( $signed( tree_1795 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1800;
always @( posedge clock ) begin
tree_1800 <= ( $signed( tree_1796 ) ) - ( $signed( tree_1797 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1801;
always @( posedge clock ) begin
tree_1801 <= ( $signed( tree_886 ) ) - ( $signed( tree_1262 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1802;
always @( posedge clock ) begin
tree_1802 <= ( $signed( tree_1798 ) ) - ( $signed( tree_1799 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1803;
always @( posedge clock ) begin
tree_1803 <= ( $signed( tree_1800 ) ) + ( $signed( tree_1801 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1804;
always @( posedge clock ) begin
tree_1804 <= ( $signed( tree_1802 ) ) + ( $signed( tree_1803 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1805;
always @( posedge clock ) begin
tree_1805 <=  - ( $signed( in[90] ) ) + ( $signed( in[99] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1806;
always @( posedge clock ) begin
tree_1806 <= ( $signed( in[105] ) ) + ( $signed( in[183] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1807;
always @( posedge clock ) begin
tree_1807 <= ( $signed( tree_1805 ) ) + ( $signed( tree_1806 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1808;
always @( posedge clock ) begin
tree_1808 <= ( $signed( tree_28 ) ) + ( $signed( tree_76 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1809;
always @( posedge clock ) begin
tree_1809 <= ( $signed( tree_14 ) ) - ( $signed( tree_41 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1810;
always @( posedge clock ) begin
tree_1810 <= ( $signed( tree_382 ) ) - ( $signed( tree_374 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1811;
always @( posedge clock ) begin
tree_1811 <=  - ( $signed( tree_130 ) ) + ( $signed( tree_578 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1812;
always @( posedge clock ) begin
tree_1812 <= ( $signed( tree_194 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1813;
always @( posedge clock ) begin
tree_1813 <= ( $signed( tree_1807 ) ) - ( $signed( tree_1808 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1814;
always @( posedge clock ) begin
tree_1814 <= ( $signed( tree_1809 ) ) + ( $signed( tree_1810 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1815;
always @( posedge clock ) begin
tree_1815 <= ( $signed( tree_1811 ) ) + ( $signed( tree_1812 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1816;
always @( posedge clock ) begin
tree_1816 <= ( $signed( tree_185 ) ) - ( $signed( tree_359 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1817;
always @( posedge clock ) begin
tree_1817 <= ( $signed( tree_883 ) ) + ( $signed( tree_861 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1818;
always @( posedge clock ) begin
tree_1818 <= ( $signed( tree_729 ) ) - ( $signed( tree_614 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1819;
always @( posedge clock ) begin
tree_1819 <=  - ( $signed( tree_966 ) ) + ( $signed( tree_474 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1820;
always @( posedge clock ) begin
tree_1820 <= ( $signed( tree_1813 ) ) + ( $signed( tree_1814 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1821;
always @( posedge clock ) begin
tree_1821 <= ( $signed( tree_1815 ) ) + ( $signed( tree_1816 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1822;
always @( posedge clock ) begin
tree_1822 <=  - ( $signed( tree_1817 ) ) + ( $signed( tree_1818 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1823;
always @( posedge clock ) begin
tree_1823 <= ( $signed( tree_1819 ) ) - ( $signed( tree_458 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1824;
always @( posedge clock ) begin
tree_1824 <= ( $signed( tree_1168 ) ) + ( $signed( tree_900 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1825;
always @( posedge clock ) begin
tree_1825 <= ( $signed( tree_1090 ) ) + ( $signed( tree_1003 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1826;
always @( posedge clock ) begin
tree_1826 <= ( $signed( tree_1820 ) ) + ( $signed( tree_1821 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1827;
always @( posedge clock ) begin
tree_1827 <= ( $signed( tree_1822 ) ) + ( $signed( tree_1823 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1828;
always @( posedge clock ) begin
tree_1828 <= ( $signed( tree_1824 ) ) + ( $signed( tree_1825 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1829;
always @( posedge clock ) begin
tree_1829 <= ( $signed( tree_1826 ) ) + ( $signed( tree_1827 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1830;
always @( posedge clock ) begin
tree_1830 <= ( $signed( tree_1828 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1831;
always @( posedge clock ) begin
tree_1831 <= ( $signed( tree_1829 ) ) - ( $signed( tree_1830 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1832;
always @( posedge clock ) begin
tree_1832 <= ( $signed( in[36] ) ) + ( $signed( in[53] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1833;
always @( posedge clock ) begin
tree_1833 <= ( $signed( in[89] ) ) + ( $signed( in[94] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1834;
always @( posedge clock ) begin
tree_1834 <= ( $signed( in[176] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1835;
always @( posedge clock ) begin
tree_1835 <= ( $signed( tree_1832 ) ) + ( $signed( tree_1833 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1836;
always @( posedge clock ) begin
tree_1836 <=  - ( $signed( tree_1834 ) ) + ( $signed( tree_203 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1837;
always @( posedge clock ) begin
tree_1837 <= ( $signed( tree_530 ) ) - ( $signed( tree_517 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1838;
always @( posedge clock ) begin
tree_1838 <= ( $signed( tree_603 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1839;
always @( posedge clock ) begin
tree_1839 <= ( $signed( tree_1835 ) ) + ( $signed( tree_1836 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1840;
always @( posedge clock ) begin
tree_1840 <= ( $signed( tree_1837 ) ) - ( $signed( tree_1838 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1841;
always @( posedge clock ) begin
tree_1841 <= ( $signed( tree_553 ) ) + ( $signed( tree_558 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1842;
always @( posedge clock ) begin
tree_1842 <= ( $signed( tree_493 ) ) - ( $signed( tree_952 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1843;
always @( posedge clock ) begin
tree_1843 <=  - ( $signed( tree_651 ) ) + ( $signed( tree_370 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1844;
always @( posedge clock ) begin
tree_1844 <= ( $signed( tree_598 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1845;
always @( posedge clock ) begin
tree_1845 <= ( $signed( tree_1839 ) ) + ( $signed( tree_1840 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1846;
always @( posedge clock ) begin
tree_1846 <=  - ( $signed( tree_1841 ) ) + ( $signed( tree_1842 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1847;
always @( posedge clock ) begin
tree_1847 <= ( $signed( tree_1843 ) ) + ( $signed( tree_1844 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1848;
always @( posedge clock ) begin
tree_1848 <= ( $signed( tree_894 ) ) + ( $signed( tree_999 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1849;
always @( posedge clock ) begin
tree_1849 <= ( $signed( tree_514 ) ) + ( $signed( tree_791 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1850;
always @( posedge clock ) begin
tree_1850 <= ( $signed( tree_1845 ) ) + ( $signed( tree_1846 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1851;
always @( posedge clock ) begin
tree_1851 <= ( $signed( tree_1847 ) ) - ( $signed( tree_1848 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1852;
always @( posedge clock ) begin
tree_1852 <= ( $signed( tree_1849 ) ) + ( $signed( tree_1617 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1853;
always @( posedge clock ) begin
tree_1853 <= ( $signed( tree_1850 ) ) + ( $signed( tree_1851 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1854;
always @( posedge clock ) begin
tree_1854 <= ( $signed( tree_1852 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1855;
always @( posedge clock ) begin
tree_1855 <= ( $signed( tree_1853 ) ) - ( $signed( tree_1854 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1856;
always @( posedge clock ) begin
tree_1856 <= ( $signed( tree_20 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1857;
always @( posedge clock ) begin
tree_1857 <= ( $signed( tree_1856 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1858;
always @( posedge clock ) begin
tree_1858 <= ( $signed( tree_1857 ) ) - ( $signed( tree_1100 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1859;
always @( posedge clock ) begin
tree_1859 <= ( $signed( tree_667 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1860;
always @( posedge clock ) begin
tree_1860 <= ( $signed( tree_1859 ) ) + ( $signed( tree_1105 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1861;
always @( posedge clock ) begin
tree_1861 <= ( $signed( tree_688 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1862;
always @( posedge clock ) begin
tree_1862 <= ( $signed( tree_1861 ) ) - ( $signed( tree_1111 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1863;
always @( posedge clock ) begin
tree_1863 <= ( $signed( in[176] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1864;
always @( posedge clock ) begin
tree_1864 <= ( $signed( tree_1863 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1865;
always @( posedge clock ) begin
tree_1865 <= ( $signed( tree_1864 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1866;
always @( posedge clock ) begin
tree_1866 <= ( $signed( tree_1865 ) ) + ( $signed( tree_1114 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1867;
always @( posedge clock ) begin
tree_1867 <= ( $signed( in[107] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1868;
always @( posedge clock ) begin
tree_1868 <= ( $signed( tree_1867 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1869;
always @( posedge clock ) begin
tree_1869 <= ( $signed( tree_1868 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1870;
always @( posedge clock ) begin
tree_1870 <= ( $signed( tree_1869 ) ) - ( $signed( tree_1125 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1871;
always @( posedge clock ) begin
tree_1871 <= ( $signed( in[135] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1872;
always @( posedge clock ) begin
tree_1872 <= ( $signed( tree_1871 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1873;
always @( posedge clock ) begin
tree_1873 <= ( $signed( tree_1872 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1874;
always @( posedge clock ) begin
tree_1874 <= ( $signed( tree_1873 ) ) - ( $signed( tree_1127 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1875;
always @( posedge clock ) begin
tree_1875 <= ( $signed( tree_719 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1876;
always @( posedge clock ) begin
tree_1876 <=  - ( $signed( tree_1875 ) ) + ( $signed( tree_1133 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1877;
always @( posedge clock ) begin
tree_1877 <= ( $signed( tree_82 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1878;
always @( posedge clock ) begin
tree_1878 <= ( $signed( tree_1877 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1879;
always @( posedge clock ) begin
tree_1879 <= ( $signed( tree_1878 ) ) + ( $signed( tree_1138 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1880;
always @( posedge clock ) begin
tree_1880 <= ( $signed( tree_742 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1881;
always @( posedge clock ) begin
tree_1881 <= ( $signed( tree_1880 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1882;
always @( posedge clock ) begin
tree_1882 <= ( $signed( tree_1881 ) ) + ( $signed( tree_1148 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1883;
always @( posedge clock ) begin
tree_1883 <= ( $signed( in[9] ) ) + ( $signed( in[20] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1884;
always @( posedge clock ) begin
tree_1884 <= ( $signed( in[74] ) ) + ( $signed( in[103] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1885;
always @( posedge clock ) begin
tree_1885 <= ( $signed( in[113] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1886;
always @( posedge clock ) begin
tree_1886 <= ( $signed( tree_1883 ) ) + ( $signed( tree_1884 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1887;
always @( posedge clock ) begin
tree_1887 <= ( $signed( tree_1885 ) ) + ( $signed( tree_76 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1888;
always @( posedge clock ) begin
tree_1888 <= ( $signed( tree_74 ) ) + ( $signed( tree_108 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1889;
always @( posedge clock ) begin
tree_1889 <= ( $signed( tree_109 ) ) - ( $signed( tree_112 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1890;
always @( posedge clock ) begin
tree_1890 <= ( $signed( tree_114 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1891;
always @( posedge clock ) begin
tree_1891 <= ( $signed( tree_1886 ) ) + ( $signed( tree_1887 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1892;
always @( posedge clock ) begin
tree_1892 <= ( $signed( tree_1888 ) ) + ( $signed( tree_1889 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1893;
always @( posedge clock ) begin
tree_1893 <= ( $signed( tree_1890 ) ) + ( $signed( tree_111 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1894;
always @( posedge clock ) begin
tree_1894 <= ( $signed( tree_746 ) ) - ( $signed( tree_749 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1895;
always @( posedge clock ) begin
tree_1895 <= ( $signed( tree_750 ) ) + ( $signed( tree_751 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1896;
always @( posedge clock ) begin
tree_1896 <= ( $signed( tree_1891 ) ) + ( $signed( tree_1892 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1897;
always @( posedge clock ) begin
tree_1897 <=  - ( $signed( tree_1893 ) ) + ( $signed( tree_1894 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1898;
always @( posedge clock ) begin
tree_1898 <= ( $signed( tree_1895 ) ) + ( $signed( tree_1110 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1899;
always @( posedge clock ) begin
tree_1899 <=  - ( $signed( tree_1151 ) ) + ( $signed( tree_748 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1900;
always @( posedge clock ) begin
tree_1900 <= ( $signed( tree_1896 ) ) + ( $signed( tree_1897 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1901;
always @( posedge clock ) begin
tree_1901 <= ( $signed( tree_1898 ) ) + ( $signed( tree_1899 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1902;
always @( posedge clock ) begin
tree_1902 <= ( $signed( tree_1153 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1903;
always @( posedge clock ) begin
tree_1903 <= ( $signed( tree_1900 ) ) + ( $signed( tree_1901 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1904;
always @( posedge clock ) begin
tree_1904 <= ( $signed( tree_1902 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1905;
always @( posedge clock ) begin
tree_1905 <= ( $signed( tree_1903 ) ) - ( $signed( tree_1904 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1906;
always @( posedge clock ) begin
tree_1906 <= ( $signed( tree_81 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1907;
always @( posedge clock ) begin
tree_1907 <= ( $signed( tree_1906 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1908;
always @( posedge clock ) begin
tree_1908 <= ( $signed( tree_1907 ) ) - ( $signed( tree_1159 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1909;
always @( posedge clock ) begin
tree_1909 <= ( $signed( in[69] ) ) + ( $signed( in[115] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1910;
always @( posedge clock ) begin
tree_1910 <= ( $signed( in[117] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1911;
always @( posedge clock ) begin
tree_1911 <=  - ( $signed( tree_1909 ) ) + ( $signed( tree_1910 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1912;
always @( posedge clock ) begin
tree_1912 <= ( $signed( tree_33 ) ) + ( $signed( tree_145 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1913;
always @( posedge clock ) begin
tree_1913 <= ( $signed( tree_31 ) ) - ( $signed( tree_148 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1914;
always @( posedge clock ) begin
tree_1914 <= ( $signed( tree_133 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1915;
always @( posedge clock ) begin
tree_1915 <= ( $signed( tree_1911 ) ) - ( $signed( tree_1912 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1916;
always @( posedge clock ) begin
tree_1916 <= ( $signed( tree_1913 ) ) - ( $signed( tree_1914 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1917;
always @( posedge clock ) begin
tree_1917 <=  - ( $signed( tree_106 ) ) + ( $signed( tree_768 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1918;
always @( posedge clock ) begin
tree_1918 <= ( $signed( tree_772 ) ) + ( $signed( tree_151 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1919;
always @( posedge clock ) begin
tree_1919 <= ( $signed( tree_157 ) ) - ( $signed( tree_160 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1920;
always @( posedge clock ) begin
tree_1920 <= ( $signed( tree_786 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1921;
always @( posedge clock ) begin
tree_1921 <= ( $signed( tree_1915 ) ) + ( $signed( tree_1916 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1922;
always @( posedge clock ) begin
tree_1922 <= ( $signed( tree_1917 ) ) + ( $signed( tree_1918 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1923;
always @( posedge clock ) begin
tree_1923 <= ( $signed( tree_1919 ) ) - ( $signed( tree_1920 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1924;
always @( posedge clock ) begin
tree_1924 <= ( $signed( tree_1165 ) ) + ( $signed( tree_1168 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1925;
always @( posedge clock ) begin
tree_1925 <= ( $signed( tree_1171 ) ) - ( $signed( tree_779 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1926;
always @( posedge clock ) begin
tree_1926 <= ( $signed( tree_781 ) ) + ( $signed( tree_1177 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1927;
always @( posedge clock ) begin
tree_1927 <=  - ( $signed( tree_1178 ) ) + ( $signed( tree_791 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1928;
always @( posedge clock ) begin
tree_1928 <= ( $signed( tree_1921 ) ) + ( $signed( tree_1922 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1929;
always @( posedge clock ) begin
tree_1929 <= ( $signed( tree_1923 ) ) - ( $signed( tree_1924 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1930;
always @( posedge clock ) begin
tree_1930 <= ( $signed( tree_1925 ) ) + ( $signed( tree_1926 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1931;
always @( posedge clock ) begin
tree_1931 <= ( $signed( tree_1927 ) ) - ( $signed( tree_1174 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1932;
always @( posedge clock ) begin
tree_1932 <= ( $signed( tree_1928 ) ) + ( $signed( tree_1929 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1933;
always @( posedge clock ) begin
tree_1933 <= ( $signed( tree_1930 ) ) + ( $signed( tree_1931 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1934;
always @( posedge clock ) begin
tree_1934 <= ( $signed( tree_1932 ) ) + ( $signed( tree_1933 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1935;
always @( posedge clock ) begin
tree_1935 <= ( $signed( in[26] ) ) + ( $signed( in[27] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1936;
always @( posedge clock ) begin
tree_1936 <= ( $signed( in[35] ) ) - ( $signed( in[111] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1937;
always @( posedge clock ) begin
tree_1937 <=  - ( $signed( in[139] ) ) + ( $signed( in[148] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1938;
always @( posedge clock ) begin
tree_1938 <= ( $signed( tree_1935 ) ) + ( $signed( tree_1936 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1939;
always @( posedge clock ) begin
tree_1939 <= ( $signed( tree_1937 ) ) + ( $signed( tree_23 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1940;
always @( posedge clock ) begin
tree_1940 <=  - ( $signed( tree_168 ) ) + ( $signed( tree_169 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1941;
always @( posedge clock ) begin
tree_1941 <= ( $signed( tree_172 ) ) - ( $signed( tree_175 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1942;
always @( posedge clock ) begin
tree_1942 <= ( $signed( tree_176 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1943;
always @( posedge clock ) begin
tree_1943 <= ( $signed( tree_1938 ) ) + ( $signed( tree_1939 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1944;
always @( posedge clock ) begin
tree_1944 <= ( $signed( tree_1940 ) ) + ( $signed( tree_1941 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1945;
always @( posedge clock ) begin
tree_1945 <= ( $signed( tree_1942 ) ) - ( $signed( tree_45 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1946;
always @( posedge clock ) begin
tree_1946 <= ( $signed( tree_171 ) ) + ( $signed( tree_655 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1947;
always @( posedge clock ) begin
tree_1947 <=  - ( $signed( tree_174 ) ) + ( $signed( tree_178 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1948;
always @( posedge clock ) begin
tree_1948 <= ( $signed( tree_180 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1949;
always @( posedge clock ) begin
tree_1949 <= ( $signed( tree_1943 ) ) + ( $signed( tree_1944 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1950;
always @( posedge clock ) begin
tree_1950 <= ( $signed( tree_1945 ) ) + ( $signed( tree_1946 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1951;
always @( posedge clock ) begin
tree_1951 <= ( $signed( tree_1947 ) ) + ( $signed( tree_1948 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1952;
always @( posedge clock ) begin
tree_1952 <= ( $signed( tree_1096 ) ) - ( $signed( tree_794 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1953;
always @( posedge clock ) begin
tree_1953 <= ( $signed( tree_779 ) ) - ( $signed( tree_796 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1954;
always @( posedge clock ) begin
tree_1954 <= ( $signed( tree_1183 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1955;
always @( posedge clock ) begin
tree_1955 <= ( $signed( tree_1949 ) ) + ( $signed( tree_1950 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1956;
always @( posedge clock ) begin
tree_1956 <= ( $signed( tree_1951 ) ) + ( $signed( tree_1952 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1957;
always @( posedge clock ) begin
tree_1957 <= ( $signed( tree_1953 ) ) + ( $signed( tree_1954 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1958;
always @( posedge clock ) begin
tree_1958 <= ( $signed( tree_1182 ) ) + ( $signed( tree_1879 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1959;
always @( posedge clock ) begin
tree_1959 <= ( $signed( tree_1955 ) ) + ( $signed( tree_1956 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1960;
always @( posedge clock ) begin
tree_1960 <= ( $signed( tree_1957 ) ) + ( $signed( tree_1958 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1961;
always @( posedge clock ) begin
tree_1961 <= ( $signed( tree_1959 ) ) + ( $signed( tree_1960 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1962;
always @( posedge clock ) begin
tree_1962 <= ( $signed( in[88] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1963;
always @( posedge clock ) begin
tree_1963 <= ( $signed( tree_1962 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1964;
always @( posedge clock ) begin
tree_1964 <= ( $signed( tree_1963 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1965;
always @( posedge clock ) begin
tree_1965 <= ( $signed( tree_1964 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1966;
always @( posedge clock ) begin
tree_1966 <= ( $signed( tree_1965 ) ) + ( $signed( tree_1189 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1967;
always @( posedge clock ) begin
tree_1967 <=  - ( $signed( in[34] ) ) + ( $signed( in[54] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1968;
always @( posedge clock ) begin
tree_1968 <= ( $signed( in[105] ) ) - ( $signed( in[180] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1969;
always @( posedge clock ) begin
tree_1969 <= ( $signed( tree_1967 ) ) + ( $signed( tree_1968 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1970;
always @( posedge clock ) begin
tree_1970 <= ( $signed( tree_38 ) ) + ( $signed( tree_14 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1971;
always @( posedge clock ) begin
tree_1971 <= ( $signed( tree_202 ) ) + ( $signed( tree_203 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1972;
always @( posedge clock ) begin
tree_1972 <= ( $signed( tree_205 ) ) + ( $signed( tree_206 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1973;
always @( posedge clock ) begin
tree_1973 <= ( $signed( tree_209 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1974;
always @( posedge clock ) begin
tree_1974 <= ( $signed( tree_1969 ) ) - ( $signed( tree_1970 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1975;
always @( posedge clock ) begin
tree_1975 <= ( $signed( tree_1971 ) ) - ( $signed( tree_1972 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1976;
always @( posedge clock ) begin
tree_1976 <= ( $signed( tree_1973 ) ) + ( $signed( tree_86 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1977;
always @( posedge clock ) begin
tree_1977 <= ( $signed( tree_106 ) ) + ( $signed( tree_776 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1978;
always @( posedge clock ) begin
tree_1978 <=  - ( $signed( tree_815 ) ) + ( $signed( tree_821 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1979;
always @( posedge clock ) begin
tree_1979 <= ( $signed( tree_822 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1980;
always @( posedge clock ) begin
tree_1980 <= ( $signed( tree_1974 ) ) + ( $signed( tree_1975 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1981;
always @( posedge clock ) begin
tree_1981 <= ( $signed( tree_1976 ) ) + ( $signed( tree_1977 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1982;
always @( posedge clock ) begin
tree_1982 <= ( $signed( tree_1978 ) ) - ( $signed( tree_1979 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1983;
always @( posedge clock ) begin
tree_1983 <= ( $signed( tree_716 ) ) + ( $signed( tree_818 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1984;
always @( posedge clock ) begin
tree_1984 <=  - ( $signed( tree_1186 ) ) + ( $signed( tree_820 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1985;
always @( posedge clock ) begin
tree_1985 <= ( $signed( tree_219 ) ) + ( $signed( tree_1102 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1986;
always @( posedge clock ) begin
tree_1986 <= ( $signed( tree_827 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1987;
always @( posedge clock ) begin
tree_1987 <= ( $signed( tree_1980 ) ) - ( $signed( tree_1981 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1988;
always @( posedge clock ) begin
tree_1988 <= ( $signed( tree_1982 ) ) - ( $signed( tree_1983 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1989;
always @( posedge clock ) begin
tree_1989 <= ( $signed( tree_1984 ) ) + ( $signed( tree_1985 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1990;
always @( posedge clock ) begin
tree_1990 <= ( $signed( tree_1986 ) ) + ( $signed( tree_1192 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1991;
always @( posedge clock ) begin
tree_1991 <= ( $signed( tree_1194 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1992;
always @( posedge clock ) begin
tree_1992 <= ( $signed( tree_1987 ) ) + ( $signed( tree_1988 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1993;
always @( posedge clock ) begin
tree_1993 <= ( $signed( tree_1989 ) ) - ( $signed( tree_1990 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1994;
always @( posedge clock ) begin
tree_1994 <= ( $signed( tree_1991 ) ) + ( $signed( tree_1198 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1995;
always @( posedge clock ) begin
tree_1995 <= ( $signed( tree_1992 ) ) + ( $signed( tree_1993 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1996;
always @( posedge clock ) begin
tree_1996 <= ( $signed( tree_1994 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_1997;
always @( posedge clock ) begin
tree_1997 <= ( $signed( tree_1995 ) ) - ( $signed( tree_1996 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1998;
always @( posedge clock ) begin
tree_1998 <=  - ( $signed( in[16] ) ) + ( $signed( in[71] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_1999;
always @( posedge clock ) begin
tree_1999 <= ( $signed( in[91] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2000;
always @( posedge clock ) begin
tree_2000 <= ( $signed( tree_1998 ) ) + ( $signed( tree_1999 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2001;
always @( posedge clock ) begin
tree_2001 <= ( $signed( tree_22 ) ) + ( $signed( tree_79 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2002;
always @( posedge clock ) begin
tree_2002 <= ( $signed( tree_225 ) ) - ( $signed( tree_226 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2003;
always @( posedge clock ) begin
tree_2003 <= ( $signed( tree_193 ) ) - ( $signed( tree_8 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2004;
always @( posedge clock ) begin
tree_2004 <= ( $signed( tree_227 ) ) - ( $signed( tree_229 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2005;
always @( posedge clock ) begin
tree_2005 <= ( $signed( tree_2000 ) ) + ( $signed( tree_2001 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2006;
always @( posedge clock ) begin
tree_2006 <= ( $signed( tree_2002 ) ) + ( $signed( tree_2003 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2007;
always @( posedge clock ) begin
tree_2007 <= ( $signed( tree_2004 ) ) + ( $signed( tree_117 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2008;
always @( posedge clock ) begin
tree_2008 <= ( $signed( tree_747 ) ) + ( $signed( tree_834 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2009;
always @( posedge clock ) begin
tree_2009 <= ( $signed( tree_235 ) ) + ( $signed( tree_50 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2010;
always @( posedge clock ) begin
tree_2010 <= ( $signed( tree_837 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2011;
always @( posedge clock ) begin
tree_2011 <= ( $signed( tree_2005 ) ) + ( $signed( tree_2006 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2012;
always @( posedge clock ) begin
tree_2012 <= ( $signed( tree_2007 ) ) + ( $signed( tree_2008 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2013;
always @( posedge clock ) begin
tree_2013 <= ( $signed( tree_2009 ) ) + ( $signed( tree_2010 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2014;
always @( posedge clock ) begin
tree_2014 <= ( $signed( tree_1199 ) ) - ( $signed( tree_1202 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2015;
always @( posedge clock ) begin
tree_2015 <= ( $signed( tree_832 ) ) - ( $signed( tree_839 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2016;
always @( posedge clock ) begin
tree_2016 <= ( $signed( tree_243 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2017;
always @( posedge clock ) begin
tree_2017 <= ( $signed( tree_2011 ) ) + ( $signed( tree_2012 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2018;
always @( posedge clock ) begin
tree_2018 <= ( $signed( tree_2013 ) ) + ( $signed( tree_2014 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2019;
always @( posedge clock ) begin
tree_2019 <= ( $signed( tree_2015 ) ) + ( $signed( tree_2016 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2020;
always @( posedge clock ) begin
tree_2020 <= ( $signed( tree_1206 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2021;
always @( posedge clock ) begin
tree_2021 <= ( $signed( tree_2017 ) ) + ( $signed( tree_2018 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2022;
always @( posedge clock ) begin
tree_2022 <= ( $signed( tree_2019 ) ) + ( $signed( tree_2020 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2023;
always @( posedge clock ) begin
tree_2023 <= ( $signed( tree_1209 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2024;
always @( posedge clock ) begin
tree_2024 <= ( $signed( tree_2021 ) ) + ( $signed( tree_2022 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2025;
always @( posedge clock ) begin
tree_2025 <= ( $signed( tree_2023 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2026;
always @( posedge clock ) begin
tree_2026 <= ( $signed( tree_2024 ) ) + ( $signed( tree_2025 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2027;
always @( posedge clock ) begin
tree_2027 <= ( $signed( tree_263 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2028;
always @( posedge clock ) begin
tree_2028 <= ( $signed( tree_2027 ) ) + ( $signed( tree_1215 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2029;
always @( posedge clock ) begin
tree_2029 <= ( $signed( tree_278 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2030;
always @( posedge clock ) begin
tree_2030 <= ( $signed( tree_2029 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2031;
always @( posedge clock ) begin
tree_2031 <= ( $signed( tree_2030 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2032;
always @( posedge clock ) begin
tree_2032 <= ( $signed( tree_2031 ) ) + ( $signed( tree_1221 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2033;
always @( posedge clock ) begin
tree_2033 <= ( $signed( tree_323 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2034;
always @( posedge clock ) begin
tree_2034 <= ( $signed( tree_2033 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2035;
always @( posedge clock ) begin
tree_2035 <=  - ( $signed( tree_2034 ) ) + ( $signed( tree_1260 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2036;
always @( posedge clock ) begin
tree_2036 <=  - ( $signed( in[62] ) ) + ( $signed( in[73] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2037;
always @( posedge clock ) begin
tree_2037 <= ( $signed( in[78] ) ) - ( $signed( in[113] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2038;
always @( posedge clock ) begin
tree_2038 <= ( $signed( in[146] ) ) + ( $signed( in[159] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2039;
always @( posedge clock ) begin
tree_2039 <= ( $signed( tree_2036 ) ) + ( $signed( tree_2037 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2040;
always @( posedge clock ) begin
tree_2040 <= ( $signed( tree_2038 ) ) + ( $signed( tree_87 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2041;
always @( posedge clock ) begin
tree_2041 <= ( $signed( tree_153 ) ) + ( $signed( tree_326 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2042;
always @( posedge clock ) begin
tree_2042 <= ( $signed( tree_327 ) ) + ( $signed( tree_328 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2043;
always @( posedge clock ) begin
tree_2043 <= ( $signed( tree_329 ) ) + ( $signed( tree_332 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2044;
always @( posedge clock ) begin
tree_2044 <= ( $signed( tree_333 ) ) + ( $signed( tree_334 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2045;
always @( posedge clock ) begin
tree_2045 <= ( $signed( tree_2039 ) ) - ( $signed( tree_2040 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2046;
always @( posedge clock ) begin
tree_2046 <= ( $signed( tree_2041 ) ) + ( $signed( tree_2042 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2047;
always @( posedge clock ) begin
tree_2047 <= ( $signed( tree_2043 ) ) - ( $signed( tree_2044 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2048;
always @( posedge clock ) begin
tree_2048 <= ( $signed( tree_712 ) ) + ( $signed( tree_672 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2049;
always @( posedge clock ) begin
tree_2049 <= ( $signed( tree_155 ) ) + ( $signed( tree_887 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2050;
always @( posedge clock ) begin
tree_2050 <= ( $signed( tree_772 ) ) + ( $signed( tree_338 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2051;
always @( posedge clock ) begin
tree_2051 <= ( $signed( tree_2045 ) ) + ( $signed( tree_2046 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2052;
always @( posedge clock ) begin
tree_2052 <= ( $signed( tree_2047 ) ) - ( $signed( tree_2048 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2053;
always @( posedge clock ) begin
tree_2053 <= ( $signed( tree_2049 ) ) - ( $signed( tree_2050 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2054;
always @( posedge clock ) begin
tree_2054 <= ( $signed( tree_890 ) ) + ( $signed( tree_1161 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2055;
always @( posedge clock ) begin
tree_2055 <=  - ( $signed( tree_872 ) ) + ( $signed( tree_856 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2056;
always @( posedge clock ) begin
tree_2056 <= ( $signed( tree_892 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2057;
always @( posedge clock ) begin
tree_2057 <= ( $signed( tree_2051 ) ) + ( $signed( tree_2052 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2058;
always @( posedge clock ) begin
tree_2058 <= ( $signed( tree_2053 ) ) + ( $signed( tree_2054 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2059;
always @( posedge clock ) begin
tree_2059 <= ( $signed( tree_2055 ) ) + ( $signed( tree_2056 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2060;
always @( posedge clock ) begin
tree_2060 <=  - ( $signed( tree_1858 ) ) + ( $signed( tree_1262 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2061;
always @( posedge clock ) begin
tree_2061 <= ( $signed( tree_2057 ) ) + ( $signed( tree_2058 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2062;
always @( posedge clock ) begin
tree_2062 <= ( $signed( tree_2059 ) ) + ( $signed( tree_2060 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2063;
always @( posedge clock ) begin
tree_2063 <= ( $signed( tree_2061 ) ) + ( $signed( tree_2062 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2064;
always @( posedge clock ) begin
tree_2064 <= ( $signed( in[0] ) ) + ( $signed( in[54] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2065;
always @( posedge clock ) begin
tree_2065 <= ( $signed( in[121] ) ) - ( $signed( in[159] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2066;
always @( posedge clock ) begin
tree_2066 <= ( $signed( in[161] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2067;
always @( posedge clock ) begin
tree_2067 <=  - ( $signed( tree_2064 ) ) + ( $signed( tree_2065 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2068;
always @( posedge clock ) begin
tree_2068 <= ( $signed( tree_2066 ) ) - ( $signed( tree_341 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2069;
always @( posedge clock ) begin
tree_2069 <=  - ( $signed( tree_316 ) ) + ( $signed( tree_342 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2070;
always @( posedge clock ) begin
tree_2070 <= ( $signed( tree_39 ) ) + ( $signed( tree_351 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2071;
always @( posedge clock ) begin
tree_2071 <= ( $signed( tree_2067 ) ) + ( $signed( tree_2068 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2072;
always @( posedge clock ) begin
tree_2072 <= ( $signed( tree_2069 ) ) - ( $signed( tree_2070 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2073;
always @( posedge clock ) begin
tree_2073 <= ( $signed( tree_159 ) ) + ( $signed( tree_697 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2074;
always @( posedge clock ) begin
tree_2074 <= ( $signed( tree_732 ) ) + ( $signed( tree_896 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2075;
always @( posedge clock ) begin
tree_2075 <= ( $signed( tree_345 ) ) - ( $signed( tree_347 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2076;
always @( posedge clock ) begin
tree_2076 <= ( $signed( tree_318 ) ) - ( $signed( tree_734 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2077;
always @( posedge clock ) begin
tree_2077 <= ( $signed( tree_656 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2078;
always @( posedge clock ) begin
tree_2078 <= ( $signed( tree_2071 ) ) + ( $signed( tree_2072 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2079;
always @( posedge clock ) begin
tree_2079 <= ( $signed( tree_2073 ) ) + ( $signed( tree_2074 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2080;
always @( posedge clock ) begin
tree_2080 <= ( $signed( tree_2075 ) ) + ( $signed( tree_2076 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2081;
always @( posedge clock ) begin
tree_2081 <=  - ( $signed( tree_2077 ) ) + ( $signed( tree_350 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2082;
always @( posedge clock ) begin
tree_2082 <= ( $signed( tree_794 ) ) + ( $signed( tree_898 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2083;
always @( posedge clock ) begin
tree_2083 <=  - ( $signed( tree_900 ) ) + ( $signed( tree_1162 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2084;
always @( posedge clock ) begin
tree_2084 <= ( $signed( tree_903 ) ) + ( $signed( tree_905 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2085;
always @( posedge clock ) begin
tree_2085 <= ( $signed( tree_1264 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2086;
always @( posedge clock ) begin
tree_2086 <= ( $signed( tree_2078 ) ) - ( $signed( tree_2079 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2087;
always @( posedge clock ) begin
tree_2087 <= ( $signed( tree_2080 ) ) + ( $signed( tree_2081 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2088;
always @( posedge clock ) begin
tree_2088 <=  - ( $signed( tree_2082 ) ) + ( $signed( tree_2083 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2089;
always @( posedge clock ) begin
tree_2089 <= ( $signed( tree_2084 ) ) + ( $signed( tree_2085 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2090;
always @( posedge clock ) begin
tree_2090 <= ( $signed( tree_2035 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2091;
always @( posedge clock ) begin
tree_2091 <= ( $signed( tree_2086 ) ) + ( $signed( tree_2087 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2092;
always @( posedge clock ) begin
tree_2092 <= ( $signed( tree_2088 ) ) - ( $signed( tree_2089 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2093;
always @( posedge clock ) begin
tree_2093 <= ( $signed( tree_2090 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2094;
always @( posedge clock ) begin
tree_2094 <= ( $signed( tree_2091 ) ) + ( $signed( tree_2092 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2095;
always @( posedge clock ) begin
tree_2095 <= ( $signed( tree_2093 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2096;
always @( posedge clock ) begin
tree_2096 <= ( $signed( tree_2094 ) ) + ( $signed( tree_2095 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2097;
always @( posedge clock ) begin
tree_2097 <= ( $signed( in[29] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2098;
always @( posedge clock ) begin
tree_2098 <= ( $signed( tree_2097 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2099;
always @( posedge clock ) begin
tree_2099 <= ( $signed( tree_2098 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2100;
always @( posedge clock ) begin
tree_2100 <= ( $signed( tree_2099 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2101;
always @( posedge clock ) begin
tree_2101 <= ( $signed( tree_2100 ) ) - ( $signed( tree_1266 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2102;
always @( posedge clock ) begin
tree_2102 <= ( $signed( in[54] ) ) + ( $signed( in[60] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2103;
always @( posedge clock ) begin
tree_2103 <= ( $signed( in[128] ) ) - ( $signed( in[135] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2104;
always @( posedge clock ) begin
tree_2104 <=  - ( $signed( in[144] ) ) + ( $signed( in[149] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2105;
always @( posedge clock ) begin
tree_2105 <= ( $signed( in[190] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2106;
always @( posedge clock ) begin
tree_2106 <= ( $signed( tree_2102 ) ) + ( $signed( tree_2103 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2107;
always @( posedge clock ) begin
tree_2107 <= ( $signed( tree_2104 ) ) - ( $signed( tree_2105 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2108;
always @( posedge clock ) begin
tree_2108 <= ( $signed( tree_74 ) ) + ( $signed( tree_18 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2109;
always @( posedge clock ) begin
tree_2109 <= ( $signed( tree_84 ) ) - ( $signed( tree_163 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2110;
always @( posedge clock ) begin
tree_2110 <= ( $signed( tree_376 ) ) - ( $signed( tree_120 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2111;
always @( posedge clock ) begin
tree_2111 <= ( $signed( tree_227 ) ) + ( $signed( tree_383 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2112;
always @( posedge clock ) begin
tree_2112 <= ( $signed( tree_2106 ) ) + ( $signed( tree_2107 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2113;
always @( posedge clock ) begin
tree_2113 <=  - ( $signed( tree_2108 ) ) + ( $signed( tree_2109 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2114;
always @( posedge clock ) begin
tree_2114 <= ( $signed( tree_2110 ) ) + ( $signed( tree_2111 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2115;
always @( posedge clock ) begin
tree_2115 <= ( $signed( tree_883 ) ) + ( $signed( tree_643 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2116;
always @( posedge clock ) begin
tree_2116 <= ( $signed( tree_377 ) ) + ( $signed( tree_379 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2117;
always @( posedge clock ) begin
tree_2117 <= ( $signed( tree_180 ) ) - ( $signed( tree_381 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2118;
always @( posedge clock ) begin
tree_2118 <= ( $signed( tree_917 ) ) + ( $signed( tree_386 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2119;
always @( posedge clock ) begin
tree_2119 <= ( $signed( tree_922 ) ) - ( $signed( tree_923 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2120;
always @( posedge clock ) begin
tree_2120 <= ( $signed( tree_2112 ) ) + ( $signed( tree_2113 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2121;
always @( posedge clock ) begin
tree_2121 <= ( $signed( tree_2114 ) ) - ( $signed( tree_2115 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2122;
always @( posedge clock ) begin
tree_2122 <=  - ( $signed( tree_2116 ) ) + ( $signed( tree_2117 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2123;
always @( posedge clock ) begin
tree_2123 <= ( $signed( tree_2118 ) ) + ( $signed( tree_2119 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2124;
always @( posedge clock ) begin
tree_2124 <= ( $signed( tree_384 ) ) + ( $signed( tree_1136 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2125;
always @( posedge clock ) begin
tree_2125 <= ( $signed( tree_2120 ) ) + ( $signed( tree_2121 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2126;
always @( posedge clock ) begin
tree_2126 <= ( $signed( tree_2122 ) ) + ( $signed( tree_2123 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2127;
always @( posedge clock ) begin
tree_2127 <=  - ( $signed( tree_2124 ) ) + ( $signed( tree_1270 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2128;
always @( posedge clock ) begin
tree_2128 <= ( $signed( tree_1272 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2129;
always @( posedge clock ) begin
tree_2129 <= ( $signed( tree_2125 ) ) + ( $signed( tree_2126 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2130;
always @( posedge clock ) begin
tree_2130 <= ( $signed( tree_2127 ) ) + ( $signed( tree_2128 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2131;
always @( posedge clock ) begin
tree_2131 <= ( $signed( tree_2032 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2132;
always @( posedge clock ) begin
tree_2132 <= ( $signed( tree_2129 ) ) + ( $signed( tree_2130 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2133;
always @( posedge clock ) begin
tree_2133 <= ( $signed( tree_2131 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2134;
always @( posedge clock ) begin
tree_2134 <= ( $signed( tree_2132 ) ) + ( $signed( tree_2133 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2135;
always @( posedge clock ) begin
tree_2135 <= ( $signed( in[51] ) ) + ( $signed( in[74] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2136;
always @( posedge clock ) begin
tree_2136 <= ( $signed( in[103] ) ) + ( $signed( in[111] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2137;
always @( posedge clock ) begin
tree_2137 <=  - ( $signed( in[121] ) ) + ( $signed( in[181] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2138;
always @( posedge clock ) begin
tree_2138 <= ( $signed( tree_2135 ) ) - ( $signed( tree_2136 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2139;
always @( posedge clock ) begin
tree_2139 <= ( $signed( tree_2137 ) ) - ( $signed( tree_153 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2140;
always @( posedge clock ) begin
tree_2140 <= ( $signed( tree_197 ) ) - ( $signed( tree_391 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2141;
always @( posedge clock ) begin
tree_2141 <= ( $signed( tree_394 ) ) - ( $signed( tree_293 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2142;
always @( posedge clock ) begin
tree_2142 <= ( $signed( tree_395 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2143;
always @( posedge clock ) begin
tree_2143 <= ( $signed( tree_2138 ) ) + ( $signed( tree_2139 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2144;
always @( posedge clock ) begin
tree_2144 <= ( $signed( tree_2140 ) ) + ( $signed( tree_2141 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2145;
always @( posedge clock ) begin
tree_2145 <= ( $signed( tree_2142 ) ) + ( $signed( tree_774 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2146;
always @( posedge clock ) begin
tree_2146 <= ( $signed( tree_36 ) ) - ( $signed( tree_678 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2147;
always @( posedge clock ) begin
tree_2147 <= ( $signed( tree_747 ) ) - ( $signed( tree_393 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2148;
always @( posedge clock ) begin
tree_2148 <= ( $signed( tree_311 ) ) + ( $signed( tree_804 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2149;
always @( posedge clock ) begin
tree_2149 <=  - ( $signed( tree_402 ) ) + ( $signed( tree_928 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2150;
always @( posedge clock ) begin
tree_2150 <= ( $signed( tree_2143 ) ) + ( $signed( tree_2144 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2151;
always @( posedge clock ) begin
tree_2151 <= ( $signed( tree_2145 ) ) + ( $signed( tree_2146 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2152;
always @( posedge clock ) begin
tree_2152 <= ( $signed( tree_2147 ) ) + ( $signed( tree_2148 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2153;
always @( posedge clock ) begin
tree_2153 <= ( $signed( tree_2149 ) ) - ( $signed( tree_1165 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2154;
always @( posedge clock ) begin
tree_2154 <=  - ( $signed( tree_368 ) ) + ( $signed( tree_925 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2155;
always @( posedge clock ) begin
tree_2155 <=  - ( $signed( tree_1274 ) ) + ( $signed( tree_399 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2156;
always @( posedge clock ) begin
tree_2156 <= ( $signed( tree_2150 ) ) + ( $signed( tree_2151 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2157;
always @( posedge clock ) begin
tree_2157 <= ( $signed( tree_2152 ) ) + ( $signed( tree_2153 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2158;
always @( posedge clock ) begin
tree_2158 <= ( $signed( tree_2154 ) ) + ( $signed( tree_2155 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2159;
always @( posedge clock ) begin
tree_2159 <= ( $signed( tree_1276 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2160;
always @( posedge clock ) begin
tree_2160 <= ( $signed( tree_2156 ) ) + ( $signed( tree_2157 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2161;
always @( posedge clock ) begin
tree_2161 <= ( $signed( tree_2158 ) ) + ( $signed( tree_2159 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2162;
always @( posedge clock ) begin
tree_2162 <= ( $signed( tree_2160 ) ) + ( $signed( tree_2161 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2163;
always @( posedge clock ) begin
tree_2163 <= ( $signed( tree_1279 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2164;
always @( posedge clock ) begin
tree_2164 <= ( $signed( tree_2162 ) ) + ( $signed( tree_2163 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2165;
always @( posedge clock ) begin
tree_2165 <= ( $signed( in[30] ) ) + ( $signed( in[56] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2166;
always @( posedge clock ) begin
tree_2166 <= ( $signed( in[163] ) ) + ( $signed( in[186] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2167;
always @( posedge clock ) begin
tree_2167 <= ( $signed( tree_2165 ) ) - ( $signed( tree_2166 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2168;
always @( posedge clock ) begin
tree_2168 <= ( $signed( tree_89 ) ) + ( $signed( tree_1 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2169;
always @( posedge clock ) begin
tree_2169 <= ( $signed( tree_41 ) ) + ( $signed( tree_225 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2170;
always @( posedge clock ) begin
tree_2170 <= ( $signed( tree_408 ) ) + ( $signed( tree_334 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2171;
always @( posedge clock ) begin
tree_2171 <= ( $signed( tree_413 ) ) + ( $signed( tree_414 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2172;
always @( posedge clock ) begin
tree_2172 <= ( $signed( tree_415 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2173;
always @( posedge clock ) begin
tree_2173 <= ( $signed( tree_2167 ) ) - ( $signed( tree_2168 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2174;
always @( posedge clock ) begin
tree_2174 <=  - ( $signed( tree_2169 ) ) + ( $signed( tree_2170 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2175;
always @( posedge clock ) begin
tree_2175 <= ( $signed( tree_2171 ) ) + ( $signed( tree_2172 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2176;
always @( posedge clock ) begin
tree_2176 <= ( $signed( tree_410 ) ) + ( $signed( tree_128 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2177;
always @( posedge clock ) begin
tree_2177 <= ( $signed( tree_753 ) ) + ( $signed( tree_936 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2178;
always @( posedge clock ) begin
tree_2178 <= ( $signed( tree_914 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2179;
always @( posedge clock ) begin
tree_2179 <= ( $signed( tree_2173 ) ) + ( $signed( tree_2174 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2180;
always @( posedge clock ) begin
tree_2180 <= ( $signed( tree_2175 ) ) + ( $signed( tree_2176 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2181;
always @( posedge clock ) begin
tree_2181 <= ( $signed( tree_2177 ) ) + ( $signed( tree_2178 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2182;
always @( posedge clock ) begin
tree_2182 <= ( $signed( tree_933 ) ) - ( $signed( tree_935 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2183;
always @( posedge clock ) begin
tree_2183 <= ( $signed( tree_820 ) ) - ( $signed( tree_939 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2184;
always @( posedge clock ) begin
tree_2184 <= ( $signed( tree_2179 ) ) + ( $signed( tree_2180 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2185;
always @( posedge clock ) begin
tree_2185 <=  - ( $signed( tree_2181 ) ) + ( $signed( tree_2182 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2186;
always @( posedge clock ) begin
tree_2186 <= ( $signed( tree_2183 ) ) + ( $signed( tree_1862 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2187;
always @( posedge clock ) begin
tree_2187 <= ( $signed( tree_1282 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2188;
always @( posedge clock ) begin
tree_2188 <= ( $signed( tree_2184 ) ) + ( $signed( tree_2185 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2189;
always @( posedge clock ) begin
tree_2189 <= ( $signed( tree_2186 ) ) + ( $signed( tree_2187 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2190;
always @( posedge clock ) begin
tree_2190 <= ( $signed( tree_2188 ) ) + ( $signed( tree_2189 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2191;
always @( posedge clock ) begin
tree_2191 <= ( $signed( in[17] ) ) - ( $signed( in[18] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2192;
always @( posedge clock ) begin
tree_2192 <= ( $signed( in[150] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2193;
always @( posedge clock ) begin
tree_2193 <= ( $signed( tree_2191 ) ) - ( $signed( tree_2192 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2194;
always @( posedge clock ) begin
tree_2194 <= ( $signed( tree_4 ) ) - ( $signed( tree_162 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2195;
always @( posedge clock ) begin
tree_2195 <=  - ( $signed( tree_99 ) ) + ( $signed( tree_122 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2196;
always @( posedge clock ) begin
tree_2196 <= ( $signed( tree_126 ) ) - ( $signed( tree_39 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2197;
always @( posedge clock ) begin
tree_2197 <= ( $signed( tree_364 ) ) + ( $signed( tree_421 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2198;
always @( posedge clock ) begin
tree_2198 <= ( $signed( tree_424 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2199;
always @( posedge clock ) begin
tree_2199 <= ( $signed( tree_2193 ) ) + ( $signed( tree_2194 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2200;
always @( posedge clock ) begin
tree_2200 <= ( $signed( tree_2195 ) ) + ( $signed( tree_2196 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2201;
always @( posedge clock ) begin
tree_2201 <= ( $signed( tree_2197 ) ) - ( $signed( tree_2198 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2202;
always @( posedge clock ) begin
tree_2202 <= ( $signed( tree_420 ) ) + ( $signed( tree_310 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2203;
always @( posedge clock ) begin
tree_2203 <= ( $signed( tree_853 ) ) + ( $signed( tree_423 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2204;
always @( posedge clock ) begin
tree_2204 <= ( $signed( tree_943 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2205;
always @( posedge clock ) begin
tree_2205 <= ( $signed( tree_2199 ) ) + ( $signed( tree_2200 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2206;
always @( posedge clock ) begin
tree_2206 <= ( $signed( tree_2201 ) ) - ( $signed( tree_2202 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2207;
always @( posedge clock ) begin
tree_2207 <= ( $signed( tree_2203 ) ) + ( $signed( tree_2204 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2208;
always @( posedge clock ) begin
tree_2208 <= ( $signed( tree_860 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2209;
always @( posedge clock ) begin
tree_2209 <= ( $signed( tree_2205 ) ) + ( $signed( tree_2206 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2210;
always @( posedge clock ) begin
tree_2210 <= ( $signed( tree_2207 ) ) + ( $signed( tree_2208 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2211;
always @( posedge clock ) begin
tree_2211 <= ( $signed( tree_1283 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2212;
always @( posedge clock ) begin
tree_2212 <= ( $signed( tree_2209 ) ) - ( $signed( tree_2210 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2213;
always @( posedge clock ) begin
tree_2213 <= ( $signed( tree_2211 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2214;
always @( posedge clock ) begin
tree_2214 <= ( $signed( tree_2212 ) ) - ( $signed( tree_2213 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2215;
always @( posedge clock ) begin
tree_2215 <= ( $signed( tree_432 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2216;
always @( posedge clock ) begin
tree_2216 <= ( $signed( tree_2215 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2217;
always @( posedge clock ) begin
tree_2217 <= ( $signed( tree_2216 ) ) - ( $signed( tree_1285 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2218;
always @( posedge clock ) begin
tree_2218 <= ( $signed( in[87] ) ) - ( $signed( in[129] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2219;
always @( posedge clock ) begin
tree_2219 <= ( $signed( tree_2218 ) ) - ( $signed( tree_152 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2220;
always @( posedge clock ) begin
tree_2220 <=  - ( $signed( tree_64 ) ) + ( $signed( tree_322 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2221;
always @( posedge clock ) begin
tree_2221 <= ( $signed( tree_17 ) ) + ( $signed( tree_126 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2222;
always @( posedge clock ) begin
tree_2222 <= ( $signed( tree_163 ) ) + ( $signed( tree_342 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2223;
always @( posedge clock ) begin
tree_2223 <= ( $signed( tree_441 ) ) + ( $signed( tree_114 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2224;
always @( posedge clock ) begin
tree_2224 <= ( $signed( tree_297 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2225;
always @( posedge clock ) begin
tree_2225 <= ( $signed( tree_2219 ) ) + ( $signed( tree_2220 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2226;
always @( posedge clock ) begin
tree_2226 <= ( $signed( tree_2221 ) ) + ( $signed( tree_2222 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2227;
always @( posedge clock ) begin
tree_2227 <= ( $signed( tree_2223 ) ) - ( $signed( tree_2224 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2228;
always @( posedge clock ) begin
tree_2228 <=  - ( $signed( tree_742 ) ) + ( $signed( tree_952 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2229;
always @( posedge clock ) begin
tree_2229 <= ( $signed( tree_440 ) ) + ( $signed( tree_850 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2230;
always @( posedge clock ) begin
tree_2230 <= ( $signed( tree_68 ) ) - ( $signed( tree_283 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2231;
always @( posedge clock ) begin
tree_2231 <= ( $signed( tree_809 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2232;
always @( posedge clock ) begin
tree_2232 <= ( $signed( tree_2225 ) ) + ( $signed( tree_2226 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2233;
always @( posedge clock ) begin
tree_2233 <= ( $signed( tree_2227 ) ) + ( $signed( tree_2228 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2234;
always @( posedge clock ) begin
tree_2234 <=  - ( $signed( tree_2229 ) ) + ( $signed( tree_2230 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2235;
always @( posedge clock ) begin
tree_2235 <= ( $signed( tree_2231 ) ) + ( $signed( tree_955 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2236;
always @( posedge clock ) begin
tree_2236 <= ( $signed( tree_445 ) ) - ( $signed( tree_827 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2237;
always @( posedge clock ) begin
tree_2237 <= ( $signed( tree_2232 ) ) + ( $signed( tree_2233 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2238;
always @( posedge clock ) begin
tree_2238 <= ( $signed( tree_2234 ) ) + ( $signed( tree_2235 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2239;
always @( posedge clock ) begin
tree_2239 <= ( $signed( tree_2236 ) ) + ( $signed( tree_1908 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2240;
always @( posedge clock ) begin
tree_2240 <= ( $signed( tree_1296 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2241;
always @( posedge clock ) begin
tree_2241 <= ( $signed( tree_2237 ) ) + ( $signed( tree_2238 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2242;
always @( posedge clock ) begin
tree_2242 <= ( $signed( tree_2239 ) ) + ( $signed( tree_2240 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2243;
always @( posedge clock ) begin
tree_2243 <= ( $signed( tree_2241 ) ) + ( $signed( tree_2242 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2244;
always @( posedge clock ) begin
tree_2244 <= ( $signed( in[41] ) ) - ( $signed( in[44] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2245;
always @( posedge clock ) begin
tree_2245 <= ( $signed( in[52] ) ) + ( $signed( in[97] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2246;
always @( posedge clock ) begin
tree_2246 <= ( $signed( in[153] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2247;
always @( posedge clock ) begin
tree_2247 <= ( $signed( tree_2244 ) ) - ( $signed( tree_2245 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2248;
always @( posedge clock ) begin
tree_2248 <= ( $signed( tree_2246 ) ) + ( $signed( tree_89 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2249;
always @( posedge clock ) begin
tree_2249 <= ( $signed( tree_199 ) ) + ( $signed( tree_169 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2250;
always @( posedge clock ) begin
tree_2250 <=  - ( $signed( tree_228 ) ) + ( $signed( tree_62 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2251;
always @( posedge clock ) begin
tree_2251 <= ( $signed( tree_221 ) ) + ( $signed( tree_270 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2252;
always @( posedge clock ) begin
tree_2252 <= ( $signed( tree_387 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2253;
always @( posedge clock ) begin
tree_2253 <= ( $signed( tree_2247 ) ) + ( $signed( tree_2248 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2254;
always @( posedge clock ) begin
tree_2254 <= ( $signed( tree_2249 ) ) + ( $signed( tree_2250 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2255;
always @( posedge clock ) begin
tree_2255 <= ( $signed( tree_2251 ) ) + ( $signed( tree_2252 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2256;
always @( posedge clock ) begin
tree_2256 <= ( $signed( tree_669 ) ) + ( $signed( tree_447 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2257;
always @( posedge clock ) begin
tree_2257 <= ( $signed( tree_303 ) ) + ( $signed( tree_966 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2258;
always @( posedge clock ) begin
tree_2258 <=  - ( $signed( tree_821 ) ) + ( $signed( tree_450 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2259;
always @( posedge clock ) begin
tree_2259 <= ( $signed( tree_2253 ) ) + ( $signed( tree_2254 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2260;
always @( posedge clock ) begin
tree_2260 <= ( $signed( tree_2255 ) ) + ( $signed( tree_2256 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2261;
always @( posedge clock ) begin
tree_2261 <= ( $signed( tree_2257 ) ) + ( $signed( tree_2258 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2262;
always @( posedge clock ) begin
tree_2262 <= ( $signed( tree_909 ) ) - ( $signed( tree_1159 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2263;
always @( posedge clock ) begin
tree_2263 <= ( $signed( tree_960 ) ) + ( $signed( tree_970 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2264;
always @( posedge clock ) begin
tree_2264 <= ( $signed( tree_2259 ) ) + ( $signed( tree_2260 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2265;
always @( posedge clock ) begin
tree_2265 <= ( $signed( tree_2261 ) ) + ( $signed( tree_2262 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2266;
always @( posedge clock ) begin
tree_2266 <= ( $signed( tree_2263 ) ) + ( $signed( tree_1305 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2267;
always @( posedge clock ) begin
tree_2267 <= ( $signed( tree_1292 ) ) + ( $signed( tree_977 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2268;
always @( posedge clock ) begin
tree_2268 <= ( $signed( tree_2264 ) ) + ( $signed( tree_2265 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2269;
always @( posedge clock ) begin
tree_2269 <= ( $signed( tree_2266 ) ) + ( $signed( tree_2267 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2270;
always @( posedge clock ) begin
tree_2270 <=  - ( $signed( tree_1301 ) ) + ( $signed( tree_1309 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2271;
always @( posedge clock ) begin
tree_2271 <= ( $signed( tree_2268 ) ) + ( $signed( tree_2269 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2272;
always @( posedge clock ) begin
tree_2272 <= ( $signed( tree_2270 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2273;
always @( posedge clock ) begin
tree_2273 <= ( $signed( tree_2271 ) ) + ( $signed( tree_2272 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2274;
always @( posedge clock ) begin
tree_2274 <=  - ( $signed( in[21] ) ) + ( $signed( in[35] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2275;
always @( posedge clock ) begin
tree_2275 <= ( $signed( in[100] ) ) - ( $signed( in[118] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2276;
always @( posedge clock ) begin
tree_2276 <= ( $signed( in[128] ) ) - ( $signed( in[160] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2277;
always @( posedge clock ) begin
tree_2277 <= ( $signed( tree_2274 ) ) + ( $signed( tree_2275 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2278;
always @( posedge clock ) begin
tree_2278 <= ( $signed( tree_2276 ) ) - ( $signed( tree_3 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2279;
always @( posedge clock ) begin
tree_2279 <= ( $signed( tree_94 ) ) - ( $signed( tree_454 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2280;
always @( posedge clock ) begin
tree_2280 <= ( $signed( tree_328 ) ) + ( $signed( tree_108 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2281;
always @( posedge clock ) begin
tree_2281 <= ( $signed( tree_193 ) ) - ( $signed( tree_404 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2282;
always @( posedge clock ) begin
tree_2282 <= ( $signed( tree_455 ) ) + ( $signed( tree_456 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2283;
always @( posedge clock ) begin
tree_2283 <= ( $signed( tree_222 ) ) - ( $signed( tree_424 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2284;
always @( posedge clock ) begin
tree_2284 <= ( $signed( tree_2277 ) ) + ( $signed( tree_2278 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2285;
always @( posedge clock ) begin
tree_2285 <= ( $signed( tree_2279 ) ) + ( $signed( tree_2280 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2286;
always @( posedge clock ) begin
tree_2286 <= ( $signed( tree_2281 ) ) + ( $signed( tree_2282 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2287;
always @( posedge clock ) begin
tree_2287 <= ( $signed( tree_2283 ) ) + ( $signed( tree_770 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2288;
always @( posedge clock ) begin
tree_2288 <=  - ( $signed( tree_768 ) ) + ( $signed( tree_239 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2289;
always @( posedge clock ) begin
tree_2289 <= ( $signed( tree_295 ) ) - ( $signed( tree_314 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2290;
always @( posedge clock ) begin
tree_2290 <= ( $signed( tree_879 ) ) + ( $signed( tree_459 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2291;
always @( posedge clock ) begin
tree_2291 <= ( $signed( tree_460 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2292;
always @( posedge clock ) begin
tree_2292 <= ( $signed( tree_2284 ) ) + ( $signed( tree_2285 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2293;
always @( posedge clock ) begin
tree_2293 <= ( $signed( tree_2286 ) ) + ( $signed( tree_2287 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2294;
always @( posedge clock ) begin
tree_2294 <= ( $signed( tree_2288 ) ) + ( $signed( tree_2289 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2295;
always @( posedge clock ) begin
tree_2295 <= ( $signed( tree_2290 ) ) + ( $signed( tree_2291 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2296;
always @( posedge clock ) begin
tree_2296 <= ( $signed( tree_842 ) ) + ( $signed( tree_428 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2297;
always @( posedge clock ) begin
tree_2297 <= ( $signed( tree_781 ) ) + ( $signed( tree_982 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2298;
always @( posedge clock ) begin
tree_2298 <= ( $signed( tree_983 ) ) + ( $signed( tree_986 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2299;
always @( posedge clock ) begin
tree_2299 <= ( $signed( tree_2292 ) ) + ( $signed( tree_2293 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2300;
always @( posedge clock ) begin
tree_2300 <= ( $signed( tree_2294 ) ) + ( $signed( tree_2295 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2301;
always @( posedge clock ) begin
tree_2301 <=  - ( $signed( tree_2296 ) ) + ( $signed( tree_2297 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2302;
always @( posedge clock ) begin
tree_2302 <=  - ( $signed( tree_2298 ) ) + ( $signed( tree_980 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2303;
always @( posedge clock ) begin
tree_2303 <= ( $signed( tree_1313 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2304;
always @( posedge clock ) begin
tree_2304 <= ( $signed( tree_2299 ) ) + ( $signed( tree_2300 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2305;
always @( posedge clock ) begin
tree_2305 <= ( $signed( tree_2301 ) ) + ( $signed( tree_2302 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2306;
always @( posedge clock ) begin
tree_2306 <= ( $signed( tree_2303 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2307;
always @( posedge clock ) begin
tree_2307 <= ( $signed( tree_2304 ) ) + ( $signed( tree_2305 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2308;
always @( posedge clock ) begin
tree_2308 <= ( $signed( tree_2306 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2309;
always @( posedge clock ) begin
tree_2309 <= ( $signed( tree_2307 ) ) - ( $signed( tree_2308 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2310;
always @( posedge clock ) begin
tree_2310 <=  - ( $signed( in[131] ) ) + ( $signed( in[148] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2311;
always @( posedge clock ) begin
tree_2311 <= ( $signed( tree_2310 ) ) + ( $signed( tree_125 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2312;
always @( posedge clock ) begin
tree_2312 <= ( $signed( tree_403 ) ) - ( $signed( tree_466 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2313;
always @( posedge clock ) begin
tree_2313 <= ( $signed( tree_467 ) ) - ( $signed( tree_451 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2314;
always @( posedge clock ) begin
tree_2314 <=  - ( $signed( tree_469 ) ) + ( $signed( tree_66 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2315;
always @( posedge clock ) begin
tree_2315 <= ( $signed( tree_2311 ) ) + ( $signed( tree_2312 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2316;
always @( posedge clock ) begin
tree_2316 <= ( $signed( tree_2313 ) ) + ( $signed( tree_2314 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2317;
always @( posedge clock ) begin
tree_2317 <=  - ( $signed( tree_463 ) ) + ( $signed( tree_465 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2318;
always @( posedge clock ) begin
tree_2318 <= ( $signed( tree_468 ) ) + ( $signed( tree_649 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2319;
always @( posedge clock ) begin
tree_2319 <= ( $signed( tree_471 ) ) - ( $signed( tree_472 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2320;
always @( posedge clock ) begin
tree_2320 <= ( $signed( tree_473 ) ) - ( $signed( tree_474 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2321;
always @( posedge clock ) begin
tree_2321 <=  - ( $signed( tree_386 ) ) + ( $signed( tree_476 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2322;
always @( posedge clock ) begin
tree_2322 <= ( $signed( tree_2315 ) ) + ( $signed( tree_2316 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2323;
always @( posedge clock ) begin
tree_2323 <= ( $signed( tree_2317 ) ) + ( $signed( tree_2318 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2324;
always @( posedge clock ) begin
tree_2324 <= ( $signed( tree_2319 ) ) + ( $signed( tree_2320 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2325;
always @( posedge clock ) begin
tree_2325 <= ( $signed( tree_2321 ) ) - ( $signed( tree_1140 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2326;
always @( posedge clock ) begin
tree_2326 <= ( $signed( tree_987 ) ) + ( $signed( tree_695 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2327;
always @( posedge clock ) begin
tree_2327 <= ( $signed( tree_989 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2328;
always @( posedge clock ) begin
tree_2328 <= ( $signed( tree_2322 ) ) + ( $signed( tree_2323 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2329;
always @( posedge clock ) begin
tree_2329 <= ( $signed( tree_2324 ) ) + ( $signed( tree_2325 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2330;
always @( posedge clock ) begin
tree_2330 <= ( $signed( tree_2326 ) ) - ( $signed( tree_2327 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2331;
always @( posedge clock ) begin
tree_2331 <= ( $signed( tree_1870 ) ) + ( $signed( tree_1206 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2332;
always @( posedge clock ) begin
tree_2332 <= ( $signed( tree_2328 ) ) + ( $signed( tree_2329 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2333;
always @( posedge clock ) begin
tree_2333 <= ( $signed( tree_2330 ) ) + ( $signed( tree_2331 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2334;
always @( posedge clock ) begin
tree_2334 <= ( $signed( tree_2332 ) ) + ( $signed( tree_2333 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2335;
always @( posedge clock ) begin
tree_2335 <= ( $signed( in[58] ) ) - ( $signed( in[62] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2336;
always @( posedge clock ) begin
tree_2336 <= ( $signed( in[88] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2337;
always @( posedge clock ) begin
tree_2337 <= ( $signed( tree_2335 ) ) + ( $signed( tree_2336 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2338;
always @( posedge clock ) begin
tree_2338 <= ( $signed( tree_6 ) ) + ( $signed( tree_115 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2339;
always @( posedge clock ) begin
tree_2339 <=  - ( $signed( tree_65 ) ) + ( $signed( tree_490 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2340;
always @( posedge clock ) begin
tree_2340 <= ( $signed( tree_536 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2341;
always @( posedge clock ) begin
tree_2341 <= ( $signed( tree_2337 ) ) + ( $signed( tree_2338 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2342;
always @( posedge clock ) begin
tree_2342 <= ( $signed( tree_2339 ) ) - ( $signed( tree_2340 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2343;
always @( posedge clock ) begin
tree_2343 <= ( $signed( tree_671 ) ) + ( $signed( tree_770 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2344;
always @( posedge clock ) begin
tree_2344 <=  - ( $signed( tree_762 ) ) + ( $signed( tree_410 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2345;
always @( posedge clock ) begin
tree_2345 <= ( $signed( tree_828 ) ) - ( $signed( tree_483 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2346;
always @( posedge clock ) begin
tree_2346 <= ( $signed( tree_846 ) ) + ( $signed( tree_539 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2347;
always @( posedge clock ) begin
tree_2347 <= ( $signed( tree_2341 ) ) + ( $signed( tree_2342 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2348;
always @( posedge clock ) begin
tree_2348 <=  - ( $signed( tree_2343 ) ) + ( $signed( tree_2344 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2349;
always @( posedge clock ) begin
tree_2349 <= ( $signed( tree_2345 ) ) - ( $signed( tree_2346 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2350;
always @( posedge clock ) begin
tree_2350 <= ( $signed( tree_533 ) ) - ( $signed( tree_1133 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2351;
always @( posedge clock ) begin
tree_2351 <= ( $signed( tree_350 ) ) + ( $signed( tree_1034 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2352;
always @( posedge clock ) begin
tree_2352 <= ( $signed( tree_1010 ) ) + ( $signed( tree_511 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2353;
always @( posedge clock ) begin
tree_2353 <= ( $signed( tree_243 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2354;
always @( posedge clock ) begin
tree_2354 <= ( $signed( tree_2347 ) ) + ( $signed( tree_2348 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2355;
always @( posedge clock ) begin
tree_2355 <= ( $signed( tree_2349 ) ) + ( $signed( tree_2350 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2356;
always @( posedge clock ) begin
tree_2356 <= ( $signed( tree_2351 ) ) + ( $signed( tree_2352 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2357;
always @( posedge clock ) begin
tree_2357 <= ( $signed( tree_2353 ) ) + ( $signed( tree_1446 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2358;
always @( posedge clock ) begin
tree_2358 <= ( $signed( tree_1032 ) ) - ( $signed( tree_1282 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2359;
always @( posedge clock ) begin
tree_2359 <= ( $signed( tree_1272 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2360;
always @( posedge clock ) begin
tree_2360 <= ( $signed( tree_2354 ) ) + ( $signed( tree_2355 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2361;
always @( posedge clock ) begin
tree_2361 <= ( $signed( tree_2356 ) ) + ( $signed( tree_2357 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2362;
always @( posedge clock ) begin
tree_2362 <= ( $signed( tree_2358 ) ) + ( $signed( tree_2359 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2363;
always @( posedge clock ) begin
tree_2363 <= ( $signed( tree_2360 ) ) + ( $signed( tree_2361 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2364;
always @( posedge clock ) begin
tree_2364 <= ( $signed( tree_2362 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2365;
always @( posedge clock ) begin
tree_2365 <= ( $signed( tree_2363 ) ) + ( $signed( tree_2364 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2366;
always @( posedge clock ) begin
tree_2366 <= ( $signed( in[158] ) ) + ( $signed( in[169] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2367;
always @( posedge clock ) begin
tree_2367 <=  - ( $signed( tree_2366 ) ) + ( $signed( tree_186 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2368;
always @( posedge clock ) begin
tree_2368 <= ( $signed( tree_304 ) ) - ( $signed( tree_77 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2369;
always @( posedge clock ) begin
tree_2369 <= ( $signed( tree_126 ) ) + ( $signed( tree_438 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2370;
always @( posedge clock ) begin
tree_2370 <=  - ( $signed( tree_448 ) ) + ( $signed( tree_545 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2371;
always @( posedge clock ) begin
tree_2371 <= ( $signed( tree_2367 ) ) + ( $signed( tree_2368 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2372;
always @( posedge clock ) begin
tree_2372 <= ( $signed( tree_2369 ) ) + ( $signed( tree_2370 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2373;
always @( posedge clock ) begin
tree_2373 <= ( $signed( tree_336 ) ) - ( $signed( tree_124 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2374;
always @( posedge clock ) begin
tree_2374 <=  - ( $signed( tree_688 ) ) + ( $signed( tree_397 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2375;
always @( posedge clock ) begin
tree_2375 <=  - ( $signed( tree_538 ) ) + ( $signed( tree_372 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2376;
always @( posedge clock ) begin
tree_2376 <= ( $signed( tree_547 ) ) + ( $signed( tree_549 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2377;
always @( posedge clock ) begin
tree_2377 <= ( $signed( tree_157 ) ) + ( $signed( tree_749 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2378;
always @( posedge clock ) begin
tree_2378 <= ( $signed( tree_922 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2379;
always @( posedge clock ) begin
tree_2379 <= ( $signed( tree_2371 ) ) + ( $signed( tree_2372 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2380;
always @( posedge clock ) begin
tree_2380 <= ( $signed( tree_2373 ) ) + ( $signed( tree_2374 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2381;
always @( posedge clock ) begin
tree_2381 <= ( $signed( tree_2375 ) ) + ( $signed( tree_2376 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2382;
always @( posedge clock ) begin
tree_2382 <=  - ( $signed( tree_2377 ) ) + ( $signed( tree_2378 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2383;
always @( posedge clock ) begin
tree_2383 <= ( $signed( tree_1028 ) ) + ( $signed( tree_551 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2384;
always @( posedge clock ) begin
tree_2384 <= ( $signed( tree_300 ) ) - ( $signed( tree_881 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2385;
always @( posedge clock ) begin
tree_2385 <= ( $signed( tree_1037 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2386;
always @( posedge clock ) begin
tree_2386 <= ( $signed( tree_2379 ) ) + ( $signed( tree_2380 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2387;
always @( posedge clock ) begin
tree_2387 <= ( $signed( tree_2381 ) ) + ( $signed( tree_2382 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2388;
always @( posedge clock ) begin
tree_2388 <=  - ( $signed( tree_2383 ) ) + ( $signed( tree_2384 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2389;
always @( posedge clock ) begin
tree_2389 <= ( $signed( tree_2385 ) ) - ( $signed( tree_1876 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2390;
always @( posedge clock ) begin
tree_2390 <= ( $signed( tree_1145 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2391;
always @( posedge clock ) begin
tree_2391 <= ( $signed( tree_2386 ) ) + ( $signed( tree_2387 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2392;
always @( posedge clock ) begin
tree_2392 <= ( $signed( tree_2388 ) ) + ( $signed( tree_2389 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2393;
always @( posedge clock ) begin
tree_2393 <= ( $signed( tree_2390 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2394;
always @( posedge clock ) begin
tree_2394 <= ( $signed( tree_2391 ) ) + ( $signed( tree_2392 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2395;
always @( posedge clock ) begin
tree_2395 <= ( $signed( tree_2393 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2396;
always @( posedge clock ) begin
tree_2396 <= ( $signed( tree_2394 ) ) + ( $signed( tree_2395 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2397;
always @( posedge clock ) begin
tree_2397 <= ( $signed( in[77] ) ) + ( $signed( in[163] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2398;
always @( posedge clock ) begin
tree_2398 <= ( $signed( in[179] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2399;
always @( posedge clock ) begin
tree_2399 <= ( $signed( tree_2397 ) ) + ( $signed( tree_2398 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2400;
always @( posedge clock ) begin
tree_2400 <= ( $signed( tree_38 ) ) + ( $signed( tree_2 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2401;
always @( posedge clock ) begin
tree_2401 <=  - ( $signed( tree_255 ) ) + ( $signed( tree_343 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2402;
always @( posedge clock ) begin
tree_2402 <= ( $signed( tree_365 ) ) + ( $signed( tree_394 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2403;
always @( posedge clock ) begin
tree_2403 <= ( $signed( tree_437 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2404;
always @( posedge clock ) begin
tree_2404 <=  - ( $signed( tree_2399 ) ) + ( $signed( tree_2400 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2405;
always @( posedge clock ) begin
tree_2405 <= ( $signed( tree_2401 ) ) - ( $signed( tree_2402 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2406;
always @( posedge clock ) begin
tree_2406 <= ( $signed( tree_2403 ) ) + ( $signed( tree_359 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2407;
always @( posedge clock ) begin
tree_2407 <=  - ( $signed( tree_678 ) ) + ( $signed( tree_117 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2408;
always @( posedge clock ) begin
tree_2408 <=  - ( $signed( tree_102 ) ) + ( $signed( tree_558 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2409;
always @( posedge clock ) begin
tree_2409 <=  - ( $signed( tree_560 ) ) + ( $signed( tree_151 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2410;
always @( posedge clock ) begin
tree_2410 <= ( $signed( tree_539 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2411;
always @( posedge clock ) begin
tree_2411 <= ( $signed( tree_2404 ) ) + ( $signed( tree_2405 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2412;
always @( posedge clock ) begin
tree_2412 <=  - ( $signed( tree_2406 ) ) + ( $signed( tree_2407 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2413;
always @( posedge clock ) begin
tree_2413 <= ( $signed( tree_2408 ) ) + ( $signed( tree_2409 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2414;
always @( posedge clock ) begin
tree_2414 <= ( $signed( tree_2410 ) ) + ( $signed( tree_556 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2415;
always @( posedge clock ) begin
tree_2415 <= ( $signed( tree_716 ) ) + ( $signed( tree_1260 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2416;
always @( posedge clock ) begin
tree_2416 <=  - ( $signed( tree_909 ) ) + ( $signed( tree_1034 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2417;
always @( posedge clock ) begin
tree_2417 <= ( $signed( tree_982 ) ) - ( $signed( tree_1040 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2418;
always @( posedge clock ) begin
tree_2418 <= ( $signed( tree_1183 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2419;
always @( posedge clock ) begin
tree_2419 <= ( $signed( tree_2411 ) ) + ( $signed( tree_2412 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2420;
always @( posedge clock ) begin
tree_2420 <= ( $signed( tree_2413 ) ) + ( $signed( tree_2414 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2421;
always @( posedge clock ) begin
tree_2421 <=  - ( $signed( tree_2415 ) ) + ( $signed( tree_2416 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2422;
always @( posedge clock ) begin
tree_2422 <= ( $signed( tree_2417 ) ) + ( $signed( tree_2418 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2423;
always @( posedge clock ) begin
tree_2423 <= ( $signed( tree_2419 ) ) + ( $signed( tree_2420 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2424;
always @( posedge clock ) begin
tree_2424 <= ( $signed( tree_2421 ) ) + ( $signed( tree_2422 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2425;
always @( posedge clock ) begin
tree_2425 <= ( $signed( tree_1882 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2426;
always @( posedge clock ) begin
tree_2426 <= ( $signed( tree_2423 ) ) + ( $signed( tree_2424 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2427;
always @( posedge clock ) begin
tree_2427 <= ( $signed( tree_2425 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2428;
always @( posedge clock ) begin
tree_2428 <= ( $signed( tree_2426 ) ) - ( $signed( tree_2427 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2429;
always @( posedge clock ) begin
tree_2429 <= ( $signed( in[33] ) ) - ( $signed( in[43] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2430;
always @( posedge clock ) begin
tree_2430 <=  - ( $signed( in[66] ) ) + ( $signed( in[177] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2431;
always @( posedge clock ) begin
tree_2431 <=  - ( $signed( in[187] ) ) + ( $signed( in[190] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2432;
always @( posedge clock ) begin
tree_2432 <= ( $signed( tree_2429 ) ) + ( $signed( tree_2430 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2433;
always @( posedge clock ) begin
tree_2433 <= ( $signed( tree_2431 ) ) + ( $signed( tree_358 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2434;
always @( posedge clock ) begin
tree_2434 <=  - ( $signed( tree_289 ) ) + ( $signed( tree_129 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2435;
always @( posedge clock ) begin
tree_2435 <= ( $signed( tree_281 ) ) - ( $signed( tree_226 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2436;
always @( posedge clock ) begin
tree_2436 <= ( $signed( tree_414 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2437;
always @( posedge clock ) begin
tree_2437 <= ( $signed( tree_2432 ) ) + ( $signed( tree_2433 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2438;
always @( posedge clock ) begin
tree_2438 <= ( $signed( tree_2434 ) ) + ( $signed( tree_2435 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2439;
always @( posedge clock ) begin
tree_2439 <= ( $signed( tree_2436 ) ) + ( $signed( tree_259 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2440;
always @( posedge clock ) begin
tree_2440 <= ( $signed( tree_285 ) ) + ( $signed( tree_321 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2441;
always @( posedge clock ) begin
tree_2441 <= ( $signed( tree_776 ) ) + ( $signed( tree_111 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2442;
always @( posedge clock ) begin
tree_2442 <=  - ( $signed( tree_759 ) ) + ( $signed( tree_354 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2443;
always @( posedge clock ) begin
tree_2443 <= ( $signed( tree_471 ) ) + ( $signed( tree_70 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2444;
always @( posedge clock ) begin
tree_2444 <= ( $signed( tree_575 ) ) + ( $signed( tree_579 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2445;
always @( posedge clock ) begin
tree_2445 <= ( $signed( tree_2437 ) ) + ( $signed( tree_2438 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2446;
always @( posedge clock ) begin
tree_2446 <=  - ( $signed( tree_2439 ) ) + ( $signed( tree_2440 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2447;
always @( posedge clock ) begin
tree_2447 <= ( $signed( tree_2441 ) ) + ( $signed( tree_2442 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2448;
always @( posedge clock ) begin
tree_2448 <= ( $signed( tree_2443 ) ) - ( $signed( tree_2444 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2449;
always @( posedge clock ) begin
tree_2449 <=  - ( $signed( tree_684 ) ) + ( $signed( tree_968 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2450;
always @( posedge clock ) begin
tree_2450 <= ( $signed( tree_574 ) ) + ( $signed( tree_1142 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2451;
always @( posedge clock ) begin
tree_2451 <=  - ( $signed( tree_1037 ) ) + ( $signed( tree_1041 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2452;
always @( posedge clock ) begin
tree_2452 <= ( $signed( tree_2445 ) ) + ( $signed( tree_2446 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2453;
always @( posedge clock ) begin
tree_2453 <= ( $signed( tree_2447 ) ) + ( $signed( tree_2448 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2454;
always @( posedge clock ) begin
tree_2454 <= ( $signed( tree_2449 ) ) + ( $signed( tree_2450 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2455;
always @( posedge clock ) begin
tree_2455 <= ( $signed( tree_2451 ) ) + ( $signed( tree_1530 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2456;
always @( posedge clock ) begin
tree_2456 <= ( $signed( tree_1043 ) ) - ( $signed( tree_1046 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2457;
always @( posedge clock ) begin
tree_2457 <= ( $signed( tree_2452 ) ) + ( $signed( tree_2453 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2458;
always @( posedge clock ) begin
tree_2458 <= ( $signed( tree_2454 ) ) + ( $signed( tree_2455 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2459;
always @( posedge clock ) begin
tree_2459 <= ( $signed( tree_2456 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2460;
always @( posedge clock ) begin
tree_2460 <= ( $signed( tree_2457 ) ) + ( $signed( tree_2458 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2461;
always @( posedge clock ) begin
tree_2461 <= ( $signed( tree_2459 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2462;
always @( posedge clock ) begin
tree_2462 <= ( $signed( tree_2460 ) ) + ( $signed( tree_2461 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2463;
always @( posedge clock ) begin
tree_2463 <= ( $signed( tree_600 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2464;
always @( posedge clock ) begin
tree_2464 <= ( $signed( tree_2463 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2465;
always @( posedge clock ) begin
tree_2465 <= ( $signed( tree_2464 ) ) + ( $signed( tree_1587 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2466;
always @( posedge clock ) begin
tree_2466 <=  - ( $signed( in[122] ) ) + ( $signed( in[178] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2467;
always @( posedge clock ) begin
tree_2467 <= ( $signed( in[182] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2468;
always @( posedge clock ) begin
tree_2468 <= ( $signed( tree_2466 ) ) - ( $signed( tree_2467 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2469;
always @( posedge clock ) begin
tree_2469 <= ( $signed( tree_76 ) ) + ( $signed( tree_14 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2470;
always @( posedge clock ) begin
tree_2470 <= ( $signed( tree_52 ) ) + ( $signed( tree_137 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2471;
always @( posedge clock ) begin
tree_2471 <= ( $signed( tree_518 ) ) + ( $signed( tree_455 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2472;
always @( posedge clock ) begin
tree_2472 <= ( $signed( tree_229 ) ) + ( $signed( tree_603 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2473;
always @( posedge clock ) begin
tree_2473 <= ( $signed( tree_481 ) ) + ( $signed( tree_383 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2474;
always @( posedge clock ) begin
tree_2474 <= ( $signed( tree_2468 ) ) - ( $signed( tree_2469 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2475;
always @( posedge clock ) begin
tree_2475 <= ( $signed( tree_2470 ) ) - ( $signed( tree_2471 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2476;
always @( posedge clock ) begin
tree_2476 <=  - ( $signed( tree_2472 ) ) + ( $signed( tree_2473 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2477;
always @( posedge clock ) begin
tree_2477 <= ( $signed( tree_447 ) ) - ( $signed( tree_336 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2478;
always @( posedge clock ) begin
tree_2478 <= ( $signed( tree_128 ) ) + ( $signed( tree_174 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2479;
always @( posedge clock ) begin
tree_2479 <= ( $signed( tree_605 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2480;
always @( posedge clock ) begin
tree_2480 <= ( $signed( tree_2474 ) ) + ( $signed( tree_2475 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2481;
always @( posedge clock ) begin
tree_2481 <= ( $signed( tree_2476 ) ) + ( $signed( tree_2477 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2482;
always @( posedge clock ) begin
tree_2482 <=  - ( $signed( tree_2478 ) ) + ( $signed( tree_2479 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2483;
always @( posedge clock ) begin
tree_2483 <= ( $signed( tree_726 ) ) + ( $signed( tree_608 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2484;
always @( posedge clock ) begin
tree_2484 <=  - ( $signed( tree_1217 ) ) + ( $signed( tree_1040 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2485;
always @( posedge clock ) begin
tree_2485 <= ( $signed( tree_699 ) ) + ( $signed( tree_1018 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2486;
always @( posedge clock ) begin
tree_2486 <= ( $signed( tree_2480 ) ) + ( $signed( tree_2481 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2487;
always @( posedge clock ) begin
tree_2487 <= ( $signed( tree_2482 ) ) + ( $signed( tree_2483 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2488;
always @( posedge clock ) begin
tree_2488 <= ( $signed( tree_2484 ) ) + ( $signed( tree_2485 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2489;
always @( posedge clock ) begin
tree_2489 <= ( $signed( tree_1446 ) ) + ( $signed( tree_1289 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2490;
always @( posedge clock ) begin
tree_2490 <= ( $signed( tree_1153 ) ) + ( $signed( tree_2028 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2491;
always @( posedge clock ) begin
tree_2491 <= ( $signed( tree_2486 ) ) + ( $signed( tree_2487 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2492;
always @( posedge clock ) begin
tree_2492 <= ( $signed( tree_2488 ) ) + ( $signed( tree_2489 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2493;
always @( posedge clock ) begin
tree_2493 <= ( $signed( tree_2490 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2494;
always @( posedge clock ) begin
tree_2494 <= ( $signed( tree_2491 ) ) + ( $signed( tree_2492 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2495;
always @( posedge clock ) begin
tree_2495 <= ( $signed( tree_2493 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2496;
always @( posedge clock ) begin
tree_2496 <= ( $signed( tree_2494 ) ) - ( $signed( tree_2495 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2497;
always @( posedge clock ) begin
tree_2497 <= ( $signed( in[38] ) ) - ( $signed( in[75] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2498;
always @( posedge clock ) begin
tree_2498 <= ( $signed( in[92] ) ) + ( $signed( in[119] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2499;
always @( posedge clock ) begin
tree_2499 <= ( $signed( tree_2497 ) ) + ( $signed( tree_2498 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2500;
always @( posedge clock ) begin
tree_2500 <= ( $signed( tree_7 ) ) - ( $signed( tree_5 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2501;
always @( posedge clock ) begin
tree_2501 <= ( $signed( tree_24 ) ) - ( $signed( tree_145 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2502;
always @( posedge clock ) begin
tree_2502 <= ( $signed( tree_298 ) ) - ( $signed( tree_343 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2503;
always @( posedge clock ) begin
tree_2503 <= ( $signed( tree_112 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2504;
always @( posedge clock ) begin
tree_2504 <= ( $signed( tree_2499 ) ) + ( $signed( tree_2500 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2505;
always @( posedge clock ) begin
tree_2505 <= ( $signed( tree_2501 ) ) + ( $signed( tree_2502 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2506;
always @( posedge clock ) begin
tree_2506 <= ( $signed( tree_2503 ) ) + ( $signed( tree_185 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2507;
always @( posedge clock ) begin
tree_2507 <=  - ( $signed( tree_690 ) ) + ( $signed( tree_240 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2508;
always @( posedge clock ) begin
tree_2508 <= ( $signed( tree_497 ) ) + ( $signed( tree_468 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2509;
always @( posedge clock ) begin
tree_2509 <=  - ( $signed( tree_917 ) ) + ( $signed( tree_612 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2510;
always @( posedge clock ) begin
tree_2510 <= ( $signed( tree_2504 ) ) + ( $signed( tree_2505 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2511;
always @( posedge clock ) begin
tree_2511 <= ( $signed( tree_2506 ) ) + ( $signed( tree_2507 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2512;
always @( posedge clock ) begin
tree_2512 <= ( $signed( tree_2508 ) ) + ( $signed( tree_2509 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2513;
always @( posedge clock ) begin
tree_2513 <= ( $signed( tree_533 ) ) + ( $signed( tree_527 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2514;
always @( posedge clock ) begin
tree_2514 <= ( $signed( tree_581 ) ) - ( $signed( tree_611 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2515;
always @( posedge clock ) begin
tree_2515 <= ( $signed( tree_898 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2516;
always @( posedge clock ) begin
tree_2516 <= ( $signed( tree_2510 ) ) + ( $signed( tree_2511 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2517;
always @( posedge clock ) begin
tree_2517 <= ( $signed( tree_2512 ) ) + ( $signed( tree_2513 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2518;
always @( posedge clock ) begin
tree_2518 <= ( $signed( tree_2514 ) ) - ( $signed( tree_2515 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2519;
always @( posedge clock ) begin
tree_2519 <= ( $signed( tree_1617 ) ) + ( $signed( tree_1296 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2520;
always @( posedge clock ) begin
tree_2520 <= ( $signed( tree_2516 ) ) + ( $signed( tree_2517 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2521;
always @( posedge clock ) begin
tree_2521 <= ( $signed( tree_2518 ) ) + ( $signed( tree_2519 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2522;
always @( posedge clock ) begin
tree_2522 <= ( $signed( tree_2520 ) ) + ( $signed( tree_2521 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2523;
always @( posedge clock ) begin
tree_2523 <= ( $signed( tree_1279 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2524;
always @( posedge clock ) begin
tree_2524 <= ( $signed( tree_2522 ) ) + ( $signed( tree_2523 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2525;
always @( posedge clock ) begin
tree_2525 <= ( $signed( in[42] ) ) + ( $signed( in[75] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2526;
always @( posedge clock ) begin
tree_2526 <= ( $signed( in[94] ) ) + ( $signed( in[140] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2527;
always @( posedge clock ) begin
tree_2527 <= ( $signed( in[170] ) ) + ( $signed( in[188] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2528;
always @( posedge clock ) begin
tree_2528 <= ( $signed( tree_2525 ) ) + ( $signed( tree_2526 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2529;
always @( posedge clock ) begin
tree_2529 <= ( $signed( tree_2527 ) ) + ( $signed( tree_57 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2530;
always @( posedge clock ) begin
tree_2530 <= ( $signed( tree_319 ) ) + ( $signed( tree_62 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2531;
always @( posedge clock ) begin
tree_2531 <= ( $signed( tree_100 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2532;
always @( posedge clock ) begin
tree_2532 <= ( $signed( tree_2528 ) ) + ( $signed( tree_2529 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2533;
always @( posedge clock ) begin
tree_2533 <= ( $signed( tree_2530 ) ) - ( $signed( tree_2531 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2534;
always @( posedge clock ) begin
tree_2534 <= ( $signed( tree_731 ) ) + ( $signed( tree_261 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2535;
always @( posedge clock ) begin
tree_2535 <= ( $signed( tree_762 ) ) + ( $signed( tree_747 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2536;
always @( posedge clock ) begin
tree_2536 <= ( $signed( tree_815 ) ) + ( $signed( tree_443 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2537;
always @( posedge clock ) begin
tree_2537 <= ( $signed( tree_614 ) ) - ( $signed( tree_509 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2538;
always @( posedge clock ) begin
tree_2538 <= ( $signed( tree_616 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2539;
always @( posedge clock ) begin
tree_2539 <= ( $signed( tree_2532 ) ) + ( $signed( tree_2533 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2540;
always @( posedge clock ) begin
tree_2540 <= ( $signed( tree_2534 ) ) + ( $signed( tree_2535 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2541;
always @( posedge clock ) begin
tree_2541 <= ( $signed( tree_2536 ) ) + ( $signed( tree_2537 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2542;
always @( posedge clock ) begin
tree_2542 <= ( $signed( tree_2538 ) ) + ( $signed( tree_428 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2543;
always @( posedge clock ) begin
tree_2543 <= ( $signed( tree_1049 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2544;
always @( posedge clock ) begin
tree_2544 <= ( $signed( tree_2539 ) ) + ( $signed( tree_2540 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2545;
always @( posedge clock ) begin
tree_2545 <= ( $signed( tree_2541 ) ) + ( $signed( tree_2542 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2546;
always @( posedge clock ) begin
tree_2546 <= ( $signed( tree_2543 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2547;
always @( posedge clock ) begin
tree_2547 <= ( $signed( tree_2544 ) ) + ( $signed( tree_2545 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2548;
always @( posedge clock ) begin
tree_2548 <= ( $signed( tree_2546 ) ) + ( $signed( tree_1966 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2549;
always @( posedge clock ) begin
tree_2549 <= ( $signed( tree_1058 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2550;
always @( posedge clock ) begin
tree_2550 <= ( $signed( tree_2547 ) ) - ( $signed( tree_2548 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2551;
always @( posedge clock ) begin
tree_2551 <= ( $signed( tree_2549 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2552;
always @( posedge clock ) begin
tree_2552 <= ( $signed( tree_2550 ) ) + ( $signed( tree_2551 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2553;
always @( posedge clock ) begin
tree_2553 <= ( $signed( in[58] ) ) + ( $signed( in[129] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2554;
always @( posedge clock ) begin
tree_2554 <= ( $signed( in[138] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2555;
always @( posedge clock ) begin
tree_2555 <=  - ( $signed( tree_2553 ) ) + ( $signed( tree_2554 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2556;
always @( posedge clock ) begin
tree_2556 <= ( $signed( tree_93 ) ) + ( $signed( tree_1 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2557;
always @( posedge clock ) begin
tree_2557 <= ( $signed( tree_382 ) ) + ( $signed( tree_175 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2558;
always @( posedge clock ) begin
tree_2558 <= ( $signed( tree_148 ) ) + ( $signed( tree_618 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2559;
always @( posedge clock ) begin
tree_2559 <= ( $signed( tree_315 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2560;
always @( posedge clock ) begin
tree_2560 <= ( $signed( tree_2555 ) ) - ( $signed( tree_2556 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2561;
always @( posedge clock ) begin
tree_2561 <= ( $signed( tree_2557 ) ) + ( $signed( tree_2558 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2562;
always @( posedge clock ) begin
tree_2562 <= ( $signed( tree_2559 ) ) + ( $signed( tree_758 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2563;
always @( posedge clock ) begin
tree_2563 <= ( $signed( tree_549 ) ) + ( $signed( tree_253 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2564;
always @( posedge clock ) begin
tree_2564 <= ( $signed( tree_928 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2565;
always @( posedge clock ) begin
tree_2565 <= ( $signed( tree_2560 ) ) - ( $signed( tree_2561 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2566;
always @( posedge clock ) begin
tree_2566 <= ( $signed( tree_2562 ) ) + ( $signed( tree_2563 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2567;
always @( posedge clock ) begin
tree_2567 <= ( $signed( tree_2564 ) ) + ( $signed( tree_710 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2568;
always @( posedge clock ) begin
tree_2568 <= ( $signed( tree_1004 ) ) + ( $signed( tree_1086 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2569;
always @( posedge clock ) begin
tree_2569 <= ( $signed( tree_2565 ) ) - ( $signed( tree_2566 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2570;
always @( posedge clock ) begin
tree_2570 <= ( $signed( tree_2567 ) ) - ( $signed( tree_2568 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2571;
always @( posedge clock ) begin
tree_2571 <= ( $signed( tree_1313 ) ) + ( $signed( tree_1088 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2572;
always @( posedge clock ) begin
tree_2572 <= ( $signed( tree_2569 ) ) + ( $signed( tree_2570 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2573;
always @( posedge clock ) begin
tree_2573 <= ( $signed( tree_2571 ) ) + ( $signed( tree_2465 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2574;
always @( posedge clock ) begin
tree_2574 <= ( $signed( tree_2572 ) ) - ( $signed( tree_2573 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2575;
always @( posedge clock ) begin
tree_2575 <= ( $signed( in[100] ) ) + ( $signed( in[114] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2576;
always @( posedge clock ) begin
tree_2576 <=  - ( $signed( in[157] ) ) + ( $signed( in[190] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2577;
always @( posedge clock ) begin
tree_2577 <= ( $signed( tree_2575 ) ) + ( $signed( tree_2576 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2578;
always @( posedge clock ) begin
tree_2578 <= ( $signed( tree_24 ) ) + ( $signed( tree_490 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2579;
always @( posedge clock ) begin
tree_2579 <=  - ( $signed( tree_270 ) ) + ( $signed( tree_617 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2580;
always @( posedge clock ) begin
tree_2580 <= ( $signed( tree_334 ) ) + ( $signed( tree_364 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2581;
always @( posedge clock ) begin
tree_2581 <= ( $signed( tree_2577 ) ) + ( $signed( tree_2578 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2582;
always @( posedge clock ) begin
tree_2582 <= ( $signed( tree_2579 ) ) + ( $signed( tree_2580 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2583;
always @( posedge clock ) begin
tree_2583 <=  - ( $signed( tree_274 ) ) + ( $signed( tree_412 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2584;
always @( posedge clock ) begin
tree_2584 <= ( $signed( tree_721 ) ) + ( $signed( tree_676 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2585;
always @( posedge clock ) begin
tree_2585 <= ( $signed( tree_729 ) ) + ( $signed( tree_541 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2586;
always @( posedge clock ) begin
tree_2586 <= ( $signed( tree_402 ) ) - ( $signed( tree_1025 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2587;
always @( posedge clock ) begin
tree_2587 <= ( $signed( tree_2581 ) ) + ( $signed( tree_2582 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2588;
always @( posedge clock ) begin
tree_2588 <= ( $signed( tree_2583 ) ) + ( $signed( tree_2584 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2589;
always @( posedge clock ) begin
tree_2589 <= ( $signed( tree_2585 ) ) + ( $signed( tree_2586 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2590;
always @( posedge clock ) begin
tree_2590 <= ( $signed( tree_551 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2591;
always @( posedge clock ) begin
tree_2591 <= ( $signed( tree_2587 ) ) + ( $signed( tree_2588 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2592;
always @( posedge clock ) begin
tree_2592 <= ( $signed( tree_2589 ) ) + ( $signed( tree_2590 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2593;
always @( posedge clock ) begin
tree_2593 <= ( $signed( tree_1192 ) ) + ( $signed( tree_592 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2594;
always @( posedge clock ) begin
tree_2594 <= ( $signed( tree_2591 ) ) + ( $signed( tree_2592 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2595;
always @( posedge clock ) begin
tree_2595 <= ( $signed( tree_2593 ) ) + ( $signed( tree_2217 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2596;
always @( posedge clock ) begin
tree_2596 <= ( $signed( tree_1309 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2597;
always @( posedge clock ) begin
tree_2597 <= ( $signed( tree_2594 ) ) + ( $signed( tree_2595 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2598;
always @( posedge clock ) begin
tree_2598 <= ( $signed( tree_2596 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2599;
always @( posedge clock ) begin
tree_2599 <= ( $signed( tree_2597 ) ) + ( $signed( tree_2598 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2600;
always @( posedge clock ) begin
tree_2600 <= ( $signed( in[2] ) ) + ( $signed( in[8] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2601;
always @( posedge clock ) begin
tree_2601 <= ( $signed( in[25] ) ) - ( $signed( in[140] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2602;
always @( posedge clock ) begin
tree_2602 <= ( $signed( in[162] ) ) - ( $signed( in[169] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2603;
always @( posedge clock ) begin
tree_2603 <= ( $signed( tree_2600 ) ) + ( $signed( tree_2601 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2604;
always @( posedge clock ) begin
tree_2604 <= ( $signed( tree_2602 ) ) + ( $signed( tree_216 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2605;
always @( posedge clock ) begin
tree_2605 <= ( $signed( tree_83 ) ) + ( $signed( tree_264 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2606;
always @( posedge clock ) begin
tree_2606 <= ( $signed( tree_601 ) ) + ( $signed( tree_149 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2607;
always @( posedge clock ) begin
tree_2607 <= ( $signed( tree_394 ) ) + ( $signed( tree_293 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2608;
always @( posedge clock ) begin
tree_2608 <=  - ( $signed( tree_545 ) ) + ( $signed( tree_250 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2609;
always @( posedge clock ) begin
tree_2609 <=  - ( $signed( tree_209 ) ) + ( $signed( tree_489 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2610;
always @( posedge clock ) begin
tree_2610 <= ( $signed( tree_2603 ) ) + ( $signed( tree_2604 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2611;
always @( posedge clock ) begin
tree_2611 <= ( $signed( tree_2605 ) ) + ( $signed( tree_2606 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2612;
always @( posedge clock ) begin
tree_2612 <= ( $signed( tree_2607 ) ) + ( $signed( tree_2608 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2613;
always @( posedge clock ) begin
tree_2613 <= ( $signed( tree_2609 ) ) + ( $signed( tree_493 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2614;
always @( posedge clock ) begin
tree_2614 <= ( $signed( tree_605 ) ) + ( $signed( tree_686 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2615;
always @( posedge clock ) begin
tree_2615 <= ( $signed( tree_473 ) ) + ( $signed( tree_1008 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2616;
always @( posedge clock ) begin
tree_2616 <= ( $signed( tree_2610 ) ) + ( $signed( tree_2611 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2617;
always @( posedge clock ) begin
tree_2617 <= ( $signed( tree_2612 ) ) + ( $signed( tree_2613 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2618;
always @( posedge clock ) begin
tree_2618 <= ( $signed( tree_2614 ) ) + ( $signed( tree_2615 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2619;
always @( posedge clock ) begin
tree_2619 <= ( $signed( tree_1090 ) ) - ( $signed( tree_1086 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2620;
always @( posedge clock ) begin
tree_2620 <= ( $signed( tree_637 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2621;
always @( posedge clock ) begin
tree_2621 <= ( $signed( tree_2616 ) ) + ( $signed( tree_2617 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2622;
always @( posedge clock ) begin
tree_2622 <= ( $signed( tree_2618 ) ) + ( $signed( tree_2619 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2623;
always @( posedge clock ) begin
tree_2623 <= ( $signed( tree_2620 ) ) - ( $signed( tree_1874 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2624;
always @( posedge clock ) begin
tree_2624 <=  - ( $signed( tree_1446 ) ) + ( $signed( tree_1046 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2625;
always @( posedge clock ) begin
tree_2625 <= ( $signed( tree_1305 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2626;
always @( posedge clock ) begin
tree_2626 <= ( $signed( tree_2621 ) ) + ( $signed( tree_2622 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2627;
always @( posedge clock ) begin
tree_2627 <= ( $signed( tree_2623 ) ) + ( $signed( tree_2624 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2628;
always @( posedge clock ) begin
tree_2628 <= ( $signed( tree_2625 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2629;
always @( posedge clock ) begin
tree_2629 <= ( $signed( tree_2626 ) ) + ( $signed( tree_2627 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2630;
always @( posedge clock ) begin
tree_2630 <= ( $signed( tree_2628 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2631;
always @( posedge clock ) begin
tree_2631 <= ( $signed( tree_2629 ) ) + ( $signed( tree_2630 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2632;
always @( posedge clock ) begin
tree_2632 <= ( $signed( in[30] ) ) + ( $signed( in[31] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2633;
always @( posedge clock ) begin
tree_2633 <= ( $signed( in[74] ) ) + ( $signed( in[114] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2634;
always @( posedge clock ) begin
tree_2634 <= ( $signed( in[161] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2635;
always @( posedge clock ) begin
tree_2635 <=  - ( $signed( tree_2632 ) ) + ( $signed( tree_2633 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2636;
always @( posedge clock ) begin
tree_2636 <= ( $signed( tree_2634 ) ) + ( $signed( tree_143 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2637;
always @( posedge clock ) begin
tree_2637 <= ( $signed( tree_147 ) ) + ( $signed( tree_168 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2638;
always @( posedge clock ) begin
tree_2638 <= ( $signed( tree_388 ) ) + ( $signed( tree_441 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2639;
always @( posedge clock ) begin
tree_2639 <= ( $signed( tree_2635 ) ) - ( $signed( tree_2636 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2640;
always @( posedge clock ) begin
tree_2640 <= ( $signed( tree_2637 ) ) + ( $signed( tree_2638 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2641;
always @( posedge clock ) begin
tree_2641 <=  - ( $signed( tree_724 ) ) + ( $signed( tree_887 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2642;
always @( posedge clock ) begin
tree_2642 <= ( $signed( tree_91 ) ) - ( $signed( tree_476 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2643;
always @( posedge clock ) begin
tree_2643 <= ( $signed( tree_2639 ) ) - ( $signed( tree_2640 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2644;
always @( posedge clock ) begin
tree_2644 <= ( $signed( tree_2641 ) ) + ( $signed( tree_2642 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2645;
always @( posedge clock ) begin
tree_2645 <= ( $signed( tree_740 ) ) + ( $signed( tree_581 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2646;
always @( posedge clock ) begin
tree_2646 <= ( $signed( tree_1274 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2647;
always @( posedge clock ) begin
tree_2647 <= ( $signed( tree_2643 ) ) + ( $signed( tree_2644 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2648;
always @( posedge clock ) begin
tree_2648 <=  - ( $signed( tree_2645 ) ) + ( $signed( tree_2646 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2649;
always @( posedge clock ) begin
tree_2649 <= ( $signed( tree_1194 ) ) - ( $signed( tree_1293 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2650;
always @( posedge clock ) begin
tree_2650 <= ( $signed( tree_2647 ) ) + ( $signed( tree_2648 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2651;
always @( posedge clock ) begin
tree_2651 <= ( $signed( tree_2649 ) ) - ( $signed( tree_2101 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2652;
always @( posedge clock ) begin
tree_2652 <= ( $signed( tree_2650 ) ) + ( $signed( tree_2651 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2653;
always @( posedge clock ) begin
tree_2653 <= ( $signed( in[94] ) ) + ( $signed( in[106] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2654;
always @( posedge clock ) begin
tree_2654 <= ( $signed( in[167] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2655;
always @( posedge clock ) begin
tree_2655 <= ( $signed( tree_2653 ) ) - ( $signed( tree_2654 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2656;
always @( posedge clock ) begin
tree_2656 <= ( $signed( tree_40 ) ) + ( $signed( tree_14 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2657;
always @( posedge clock ) begin
tree_2657 <= ( $signed( tree_255 ) ) + ( $signed( tree_125 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2658;
always @( posedge clock ) begin
tree_2658 <= ( $signed( tree_352 ) ) - ( $signed( tree_120 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2659;
always @( posedge clock ) begin
tree_2659 <= ( $signed( tree_51 ) ) - ( $signed( tree_491 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2660;
always @( posedge clock ) begin
tree_2660 <= ( $signed( tree_585 ) ) + ( $signed( tree_503 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2661;
always @( posedge clock ) begin
tree_2661 <= ( $signed( tree_2655 ) ) + ( $signed( tree_2656 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2662;
always @( posedge clock ) begin
tree_2662 <= ( $signed( tree_2657 ) ) + ( $signed( tree_2658 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2663;
always @( posedge clock ) begin
tree_2663 <= ( $signed( tree_2659 ) ) + ( $signed( tree_2660 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2664;
always @( posedge clock ) begin
tree_2664 <= ( $signed( tree_714 ) ) - ( $signed( tree_804 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2665;
always @( posedge clock ) begin
tree_2665 <= ( $signed( tree_178 ) ) + ( $signed( tree_596 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2666;
always @( posedge clock ) begin
tree_2666 <= ( $signed( tree_235 ) ) + ( $signed( tree_631 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2667;
always @( posedge clock ) begin
tree_2667 <= ( $signed( tree_450 ) ) - ( $signed( tree_751 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2668;
always @( posedge clock ) begin
tree_2668 <= ( $signed( tree_2661 ) ) + ( $signed( tree_2662 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2669;
always @( posedge clock ) begin
tree_2669 <= ( $signed( tree_2663 ) ) + ( $signed( tree_2664 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2670;
always @( posedge clock ) begin
tree_2670 <= ( $signed( tree_2665 ) ) + ( $signed( tree_2666 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2671;
always @( posedge clock ) begin
tree_2671 <= ( $signed( tree_2667 ) ) + ( $signed( tree_556 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2672;
always @( posedge clock ) begin
tree_2672 <= ( $signed( tree_533 ) ) + ( $signed( tree_1171 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2673;
always @( posedge clock ) begin
tree_2673 <= ( $signed( tree_735 ) ) - ( $signed( tree_983 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2674;
always @( posedge clock ) begin
tree_2674 <= ( $signed( tree_637 ) ) + ( $signed( tree_445 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2675;
always @( posedge clock ) begin
tree_2675 <= ( $signed( tree_915 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2676;
always @( posedge clock ) begin
tree_2676 <= ( $signed( tree_2668 ) ) + ( $signed( tree_2669 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2677;
always @( posedge clock ) begin
tree_2677 <= ( $signed( tree_2670 ) ) + ( $signed( tree_2671 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2678;
always @( posedge clock ) begin
tree_2678 <= ( $signed( tree_2672 ) ) + ( $signed( tree_2673 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2679;
always @( posedge clock ) begin
tree_2679 <= ( $signed( tree_2674 ) ) + ( $signed( tree_2675 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2680;
always @( posedge clock ) begin
tree_2680 <= ( $signed( tree_1866 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2681;
always @( posedge clock ) begin
tree_2681 <= ( $signed( tree_2676 ) ) + ( $signed( tree_2677 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2682;
always @( posedge clock ) begin
tree_2682 <= ( $signed( tree_2678 ) ) + ( $signed( tree_2679 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2683;
always @( posedge clock ) begin
tree_2683 <= ( $signed( tree_2680 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2684;
always @( posedge clock ) begin
tree_2684 <= ( $signed( tree_2681 ) ) + ( $signed( tree_2682 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2685;
always @( posedge clock ) begin
tree_2685 <= ( $signed( tree_2683 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2686;
always @( posedge clock ) begin
tree_2686 <= ( $signed( tree_2684 ) ) + ( $signed( tree_2685 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2687;
always @( posedge clock ) begin
tree_2687 <= ( $signed( in[136] ) ) + ( $signed( in[150] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2688;
always @( posedge clock ) begin
tree_2688 <= ( $signed( in[166] ) ) + ( $signed( in[181] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2689;
always @( posedge clock ) begin
tree_2689 <= ( $signed( tree_2687 ) ) + ( $signed( tree_2688 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2690;
always @( posedge clock ) begin
tree_2690 <= ( $signed( tree_0 ) ) - ( $signed( tree_1 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2691;
always @( posedge clock ) begin
tree_2691 <= ( $signed( tree_2 ) ) - ( $signed( tree_3 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2692;
always @( posedge clock ) begin
tree_2692 <= ( $signed( tree_8 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2693;
always @( posedge clock ) begin
tree_2693 <=  - ( $signed( tree_2689 ) ) + ( $signed( tree_2690 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2694;
always @( posedge clock ) begin
tree_2694 <= ( $signed( tree_2691 ) ) - ( $signed( tree_2692 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2695;
always @( posedge clock ) begin
tree_2695 <= ( $signed( tree_641 ) ) + ( $signed( tree_643 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2696;
always @( posedge clock ) begin
tree_2696 <= ( $signed( tree_646 ) ) + ( $signed( tree_647 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2697;
always @( posedge clock ) begin
tree_2697 <= ( $signed( tree_649 ) ) - ( $signed( tree_651 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2698;
always @( posedge clock ) begin
tree_2698 <= ( $signed( tree_653 ) ) + ( $signed( tree_656 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2699;
always @( posedge clock ) begin
tree_2699 <= ( $signed( tree_661 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2700;
always @( posedge clock ) begin
tree_2700 <= ( $signed( tree_2693 ) ) + ( $signed( tree_2694 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2701;
always @( posedge clock ) begin
tree_2701 <= ( $signed( tree_2695 ) ) + ( $signed( tree_2696 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2702;
always @( posedge clock ) begin
tree_2702 <= ( $signed( tree_2697 ) ) - ( $signed( tree_2698 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2703;
always @( posedge clock ) begin
tree_2703 <= ( $signed( tree_2699 ) ) + ( $signed( tree_1093 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2704;
always @( posedge clock ) begin
tree_2704 <=  - ( $signed( tree_1096 ) ) + ( $signed( tree_1098 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2705;
always @( posedge clock ) begin
tree_2705 <= ( $signed( tree_1102 ) ) - ( $signed( tree_1103 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2706;
always @( posedge clock ) begin
tree_2706 <= ( $signed( tree_2700 ) ) - ( $signed( tree_2701 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2707;
always @( posedge clock ) begin
tree_2707 <= ( $signed( tree_2702 ) ) - ( $signed( tree_2703 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2708;
always @( posedge clock ) begin
tree_2708 <= ( $signed( tree_2704 ) ) + ( $signed( tree_2705 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2709;
always @( posedge clock ) begin
tree_2709 <= ( $signed( tree_1858 ) ) + ( $signed( tree_1860 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2710;
always @( posedge clock ) begin
tree_2710 <= ( $signed( tree_2706 ) ) + ( $signed( tree_2707 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2711;
always @( posedge clock ) begin
tree_2711 <= ( $signed( tree_2708 ) ) - ( $signed( tree_2709 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2712;
always @( posedge clock ) begin
tree_2712 <= ( $signed( tree_2710 ) ) + ( $signed( tree_2711 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2713;
always @( posedge clock ) begin
tree_2713 <= ( $signed( in[9] ) ) + ( $signed( in[76] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2714;
always @( posedge clock ) begin
tree_2714 <= ( $signed( in[132] ) ) - ( $signed( in[191] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2715;
always @( posedge clock ) begin
tree_2715 <= ( $signed( tree_2713 ) ) + ( $signed( tree_2714 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2716;
always @( posedge clock ) begin
tree_2716 <=  - ( $signed( tree_32 ) ) + ( $signed( tree_17 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2717;
always @( posedge clock ) begin
tree_2717 <=  - ( $signed( tree_33 ) ) + ( $signed( tree_25 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2718;
always @( posedge clock ) begin
tree_2718 <= ( $signed( tree_39 ) ) + ( $signed( tree_43 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2719;
always @( posedge clock ) begin
tree_2719 <= ( $signed( tree_48 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2720;
always @( posedge clock ) begin
tree_2720 <= ( $signed( tree_2715 ) ) + ( $signed( tree_2716 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2721;
always @( posedge clock ) begin
tree_2721 <= ( $signed( tree_2717 ) ) + ( $signed( tree_2718 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2722;
always @( posedge clock ) begin
tree_2722 <=  - ( $signed( tree_2719 ) ) + ( $signed( tree_671 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2723;
always @( posedge clock ) begin
tree_2723 <= ( $signed( tree_36 ) ) - ( $signed( tree_674 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2724;
always @( posedge clock ) begin
tree_2724 <= ( $signed( tree_676 ) ) + ( $signed( tree_50 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2725;
always @( posedge clock ) begin
tree_2725 <= ( $signed( tree_686 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2726;
always @( posedge clock ) begin
tree_2726 <= ( $signed( tree_2720 ) ) + ( $signed( tree_2721 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2727;
always @( posedge clock ) begin
tree_2727 <= ( $signed( tree_2722 ) ) + ( $signed( tree_2723 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2728;
always @( posedge clock ) begin
tree_2728 <= ( $signed( tree_2724 ) ) - ( $signed( tree_2725 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2729;
always @( posedge clock ) begin
tree_2729 <= ( $signed( tree_1108 ) ) - ( $signed( tree_1110 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2730;
always @( posedge clock ) begin
tree_2730 <=  - ( $signed( tree_681 ) ) + ( $signed( tree_684 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2731;
always @( posedge clock ) begin
tree_2731 <= ( $signed( tree_695 ) ) + ( $signed( tree_699 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2732;
always @( posedge clock ) begin
tree_2732 <= ( $signed( tree_2726 ) ) + ( $signed( tree_2727 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2733;
always @( posedge clock ) begin
tree_2733 <= ( $signed( tree_2728 ) ) + ( $signed( tree_2729 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2734;
always @( posedge clock ) begin
tree_2734 <= ( $signed( tree_2730 ) ) + ( $signed( tree_2731 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2735;
always @( posedge clock ) begin
tree_2735 <= ( $signed( tree_1862 ) ) + ( $signed( tree_1866 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2736;
always @( posedge clock ) begin
tree_2736 <= ( $signed( tree_2732 ) ) + ( $signed( tree_2733 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2737;
always @( posedge clock ) begin
tree_2737 <= ( $signed( tree_2734 ) ) + ( $signed( tree_2735 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2738;
always @( posedge clock ) begin
tree_2738 <= ( $signed( tree_2736 ) ) + ( $signed( tree_2737 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2739;
always @( posedge clock ) begin
tree_2739 <= ( $signed( tree_74 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2740;
always @( posedge clock ) begin
tree_2740 <= ( $signed( tree_2739 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2741;
always @( posedge clock ) begin
tree_2741 <= ( $signed( tree_2740 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2742;
always @( posedge clock ) begin
tree_2742 <= ( $signed( tree_2741 ) ) - ( $signed( tree_1870 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2743;
always @( posedge clock ) begin
tree_2743 <= ( $signed( tree_1874 ) ) - ( $signed( tree_1130 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2744;
always @( posedge clock ) begin
tree_2744 <= ( $signed( in[28] ) ) + ( $signed( in[34] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2745;
always @( posedge clock ) begin
tree_2745 <= ( $signed( in[73] ) ) + ( $signed( in[84] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2746;
always @( posedge clock ) begin
tree_2746 <=  - ( $signed( in[173] ) ) + ( $signed( in[189] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2747;
always @( posedge clock ) begin
tree_2747 <=  - ( $signed( tree_2744 ) ) + ( $signed( tree_2745 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2748;
always @( posedge clock ) begin
tree_2748 <= ( $signed( tree_2746 ) ) + ( $signed( tree_41 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2749;
always @( posedge clock ) begin
tree_2749 <= ( $signed( tree_92 ) ) + ( $signed( tree_100 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2750;
always @( posedge clock ) begin
tree_2750 <= ( $signed( tree_2747 ) ) + ( $signed( tree_2748 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2751;
always @( posedge clock ) begin
tree_2751 <=  - ( $signed( tree_2749 ) ) + ( $signed( tree_86 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2752;
always @( posedge clock ) begin
tree_2752 <= ( $signed( tree_701 ) ) + ( $signed( tree_728 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2753;
always @( posedge clock ) begin
tree_2753 <=  - ( $signed( tree_91 ) ) + ( $signed( tree_729 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2754;
always @( posedge clock ) begin
tree_2754 <= ( $signed( tree_734 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2755;
always @( posedge clock ) begin
tree_2755 <= ( $signed( tree_2750 ) ) + ( $signed( tree_2751 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2756;
always @( posedge clock ) begin
tree_2756 <=  - ( $signed( tree_2752 ) ) + ( $signed( tree_2753 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2757;
always @( posedge clock ) begin
tree_2757 <= ( $signed( tree_2754 ) ) + ( $signed( tree_1140 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2758;
always @( posedge clock ) begin
tree_2758 <=  - ( $signed( tree_726 ) ) + ( $signed( tree_1141 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2759;
always @( posedge clock ) begin
tree_2759 <= ( $signed( tree_735 ) ) + ( $signed( tree_1142 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2760;
always @( posedge clock ) begin
tree_2760 <= ( $signed( tree_2755 ) ) + ( $signed( tree_2756 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2761;
always @( posedge clock ) begin
tree_2761 <= ( $signed( tree_2757 ) ) + ( $signed( tree_2758 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2762;
always @( posedge clock ) begin
tree_2762 <= ( $signed( tree_2759 ) ) + ( $signed( tree_1145 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2763;
always @( posedge clock ) begin
tree_2763 <= ( $signed( tree_2760 ) ) + ( $signed( tree_2761 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2764;
always @( posedge clock ) begin
tree_2764 <= ( $signed( tree_2762 ) ) + ( $signed( tree_1882 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2765;
always @( posedge clock ) begin
tree_2765 <= ( $signed( tree_2763 ) ) - ( $signed( tree_2764 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2766;
always @( posedge clock ) begin
tree_2766 <= ( $signed( in[68] ) ) + ( $signed( in[75] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2767;
always @( posedge clock ) begin
tree_2767 <=  - ( $signed( in[80] ) ) + ( $signed( in[112] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2768;
always @( posedge clock ) begin
tree_2768 <= ( $signed( tree_2766 ) ) + ( $signed( tree_2767 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2769;
always @( posedge clock ) begin
tree_2769 <= ( $signed( tree_125 ) ) + ( $signed( tree_126 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2770;
always @( posedge clock ) begin
tree_2770 <= ( $signed( tree_129 ) ) + ( $signed( tree_130 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2771;
always @( posedge clock ) begin
tree_2771 <=  - ( $signed( tree_131 ) ) + ( $signed( tree_132 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2772;
always @( posedge clock ) begin
tree_2772 <= ( $signed( tree_133 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2773;
always @( posedge clock ) begin
tree_2773 <= ( $signed( tree_2768 ) ) + ( $signed( tree_2769 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2774;
always @( posedge clock ) begin
tree_2774 <= ( $signed( tree_2770 ) ) + ( $signed( tree_2771 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2775;
always @( posedge clock ) begin
tree_2775 <= ( $signed( tree_2772 ) ) + ( $signed( tree_98 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2776;
always @( posedge clock ) begin
tree_2776 <= ( $signed( tree_128 ) ) - ( $signed( tree_757 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2777;
always @( posedge clock ) begin
tree_2777 <= ( $signed( tree_760 ) ) + ( $signed( tree_764 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2778;
always @( posedge clock ) begin
tree_2778 <= ( $signed( tree_2773 ) ) + ( $signed( tree_2774 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2779;
always @( posedge clock ) begin
tree_2779 <= ( $signed( tree_2775 ) ) + ( $signed( tree_2776 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2780;
always @( posedge clock ) begin
tree_2780 <= ( $signed( tree_2777 ) ) + ( $signed( tree_684 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2781;
always @( posedge clock ) begin
tree_2781 <= ( $signed( tree_1138 ) ) + ( $signed( tree_1161 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2782;
always @( posedge clock ) begin
tree_2782 <= ( $signed( tree_1162 ) ) - ( $signed( tree_766 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2783;
always @( posedge clock ) begin
tree_2783 <= ( $signed( tree_2778 ) ) + ( $signed( tree_2779 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2784;
always @( posedge clock ) begin
tree_2784 <= ( $signed( tree_2780 ) ) + ( $signed( tree_2781 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2785;
always @( posedge clock ) begin
tree_2785 <= ( $signed( tree_2782 ) ) + ( $signed( tree_1156 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2786;
always @( posedge clock ) begin
tree_2786 <=  - ( $signed( tree_1908 ) ) + ( $signed( tree_1860 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2787;
always @( posedge clock ) begin
tree_2787 <= ( $signed( tree_2783 ) ) + ( $signed( tree_2784 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2788;
always @( posedge clock ) begin
tree_2788 <= ( $signed( tree_2785 ) ) + ( $signed( tree_2786 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2789;
always @( posedge clock ) begin
tree_2789 <= ( $signed( tree_2787 ) ) + ( $signed( tree_2788 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2790;
always @( posedge clock ) begin
tree_2790 <= ( $signed( tree_813 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2791;
always @( posedge clock ) begin
tree_2791 <= ( $signed( tree_2790 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2792;
always @( posedge clock ) begin
tree_2792 <= ( $signed( tree_2791 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2793;
always @( posedge clock ) begin
tree_2793 <= ( $signed( tree_2792 ) ) + ( $signed( tree_1966 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2794;
always @( posedge clock ) begin
tree_2794 <=  - ( $signed( in[36] ) ) + ( $signed( in[37] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2795;
always @( posedge clock ) begin
tree_2795 <=  - ( $signed( in[113] ) ) + ( $signed( in[121] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2796;
always @( posedge clock ) begin
tree_2796 <= ( $signed( in[168] ) ) + ( $signed( in[191] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2797;
always @( posedge clock ) begin
tree_2797 <= ( $signed( tree_2794 ) ) + ( $signed( tree_2795 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2798;
always @( posedge clock ) begin
tree_2798 <=  - ( $signed( tree_2796 ) ) + ( $signed( tree_187 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2799;
always @( posedge clock ) begin
tree_2799 <= ( $signed( tree_54 ) ) + ( $signed( tree_60 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2800;
always @( posedge clock ) begin
tree_2800 <= ( $signed( tree_244 ) ) + ( $signed( tree_250 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2801;
always @( posedge clock ) begin
tree_2801 <= ( $signed( tree_251 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2802;
always @( posedge clock ) begin
tree_2802 <= ( $signed( tree_2797 ) ) + ( $signed( tree_2798 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2803;
always @( posedge clock ) begin
tree_2803 <=  - ( $signed( tree_2799 ) ) + ( $signed( tree_2800 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2804;
always @( posedge clock ) begin
tree_2804 <= ( $signed( tree_2801 ) ) + ( $signed( tree_705 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2805;
always @( posedge clock ) begin
tree_2805 <= ( $signed( tree_246 ) ) + ( $signed( tree_253 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2806;
always @( posedge clock ) begin
tree_2806 <= ( $signed( tree_846 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2807;
always @( posedge clock ) begin
tree_2807 <= ( $signed( tree_2802 ) ) + ( $signed( tree_2803 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2808;
always @( posedge clock ) begin
tree_2808 <=  - ( $signed( tree_2804 ) ) + ( $signed( tree_2805 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2809;
always @( posedge clock ) begin
tree_2809 <= ( $signed( tree_2806 ) ) + ( $signed( tree_842 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2810;
always @( posedge clock ) begin
tree_2810 <=  - ( $signed( tree_844 ) ) + ( $signed( tree_249 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2811;
always @( posedge clock ) begin
tree_2811 <= ( $signed( tree_848 ) ) + ( $signed( tree_1212 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2812;
always @( posedge clock ) begin
tree_2812 <= ( $signed( tree_2807 ) ) + ( $signed( tree_2808 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2813;
always @( posedge clock ) begin
tree_2813 <= ( $signed( tree_2809 ) ) + ( $signed( tree_2810 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2814;
always @( posedge clock ) begin
tree_2814 <=  - ( $signed( tree_2811 ) ) + ( $signed( tree_1870 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2815;
always @( posedge clock ) begin
tree_2815 <= ( $signed( tree_1214 ) ) + ( $signed( tree_2028 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2816;
always @( posedge clock ) begin
tree_2816 <= ( $signed( tree_2812 ) ) + ( $signed( tree_2813 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2817;
always @( posedge clock ) begin
tree_2817 <= ( $signed( tree_2814 ) ) + ( $signed( tree_2815 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2818;
always @( posedge clock ) begin
tree_2818 <= ( $signed( tree_2816 ) ) + ( $signed( tree_2817 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2819;
always @( posedge clock ) begin
tree_2819 <= ( $signed( in[74] ) ) + ( $signed( in[174] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2820;
always @( posedge clock ) begin
tree_2820 <= ( $signed( tree_2819 ) ) - ( $signed( tree_28 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2821;
always @( posedge clock ) begin
tree_2821 <=  - ( $signed( tree_25 ) ) + ( $signed( tree_233 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2822;
always @( posedge clock ) begin
tree_2822 <= ( $signed( tree_104 ) ) + ( $signed( tree_270 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2823;
always @( posedge clock ) begin
tree_2823 <=  - ( $signed( tree_271 ) ) + ( $signed( tree_272 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2824;
always @( posedge clock ) begin
tree_2824 <= ( $signed( tree_2820 ) ) + ( $signed( tree_2821 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2825;
always @( posedge clock ) begin
tree_2825 <= ( $signed( tree_2822 ) ) + ( $signed( tree_2823 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2826;
always @( posedge clock ) begin
tree_2826 <= ( $signed( tree_267 ) ) + ( $signed( tree_269 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2827;
always @( posedge clock ) begin
tree_2827 <= ( $signed( tree_2824 ) ) + ( $signed( tree_2825 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2828;
always @( posedge clock ) begin
tree_2828 <= ( $signed( tree_2826 ) ) - ( $signed( tree_716 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2829;
always @( posedge clock ) begin
tree_2829 <= ( $signed( tree_856 ) ) + ( $signed( tree_1217 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2830;
always @( posedge clock ) begin
tree_2830 <= ( $signed( tree_860 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2831;
always @( posedge clock ) begin
tree_2831 <= ( $signed( tree_2827 ) ) + ( $signed( tree_2828 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2832;
always @( posedge clock ) begin
tree_2832 <= ( $signed( tree_2829 ) ) + ( $signed( tree_2830 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2833;
always @( posedge clock ) begin
tree_2833 <= ( $signed( tree_2831 ) ) + ( $signed( tree_2832 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2834;
always @( posedge clock ) begin
tree_2834 <= ( $signed( tree_2032 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2835;
always @( posedge clock ) begin
tree_2835 <= ( $signed( tree_2833 ) ) + ( $signed( tree_2834 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2836;
always @( posedge clock ) begin
tree_2836 <= ( $signed( in[8] ) ) - ( $signed( in[16] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2837;
always @( posedge clock ) begin
tree_2837 <= ( $signed( in[47] ) ) + ( $signed( in[65] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2838;
always @( posedge clock ) begin
tree_2838 <= ( $signed( in[77] ) ) + ( $signed( in[88] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2839;
always @( posedge clock ) begin
tree_2839 <= ( $signed( in[146] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2840;
always @( posedge clock ) begin
tree_2840 <= ( $signed( tree_2836 ) ) - ( $signed( tree_2837 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2841;
always @( posedge clock ) begin
tree_2841 <=  - ( $signed( tree_2838 ) ) + ( $signed( tree_2839 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2842;
always @( posedge clock ) begin
tree_2842 <= ( $signed( tree_30 ) ) - ( $signed( tree_29 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2843;
always @( posedge clock ) begin
tree_2843 <= ( $signed( tree_93 ) ) + ( $signed( tree_281 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2844;
always @( posedge clock ) begin
tree_2844 <= ( $signed( tree_176 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2845;
always @( posedge clock ) begin
tree_2845 <= ( $signed( tree_2840 ) ) + ( $signed( tree_2841 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2846;
always @( posedge clock ) begin
tree_2846 <= ( $signed( tree_2842 ) ) + ( $signed( tree_2843 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2847;
always @( posedge clock ) begin
tree_2847 <= ( $signed( tree_2844 ) ) + ( $signed( tree_639 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2848;
always @( posedge clock ) begin
tree_2848 <= ( $signed( tree_45 ) ) + ( $signed( tree_279 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2849;
always @( posedge clock ) begin
tree_2849 <= ( $signed( tree_861 ) ) + ( $signed( tree_753 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2850;
always @( posedge clock ) begin
tree_2850 <= ( $signed( tree_282 ) ) - ( $signed( tree_653 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2851;
always @( posedge clock ) begin
tree_2851 <= ( $signed( tree_283 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2852;
always @( posedge clock ) begin
tree_2852 <= ( $signed( tree_2845 ) ) + ( $signed( tree_2846 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2853;
always @( posedge clock ) begin
tree_2853 <= ( $signed( tree_2847 ) ) + ( $signed( tree_2848 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2854;
always @( posedge clock ) begin
tree_2854 <= ( $signed( tree_2849 ) ) + ( $signed( tree_2850 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2855;
always @( posedge clock ) begin
tree_2855 <= ( $signed( tree_2851 ) ) - ( $signed( tree_862 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2856;
always @( posedge clock ) begin
tree_2856 <= ( $signed( tree_2852 ) ) - ( $signed( tree_2853 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2857;
always @( posedge clock ) begin
tree_2857 <= ( $signed( tree_2854 ) ) + ( $signed( tree_2855 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2858;
always @( posedge clock ) begin
tree_2858 <= ( $signed( tree_1223 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2859;
always @( posedge clock ) begin
tree_2859 <= ( $signed( tree_2856 ) ) + ( $signed( tree_2857 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2860;
always @( posedge clock ) begin
tree_2860 <=  - ( $signed( tree_2858 ) ) + ( $signed( tree_2742 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2861;
always @( posedge clock ) begin
tree_2861 <= ( $signed( tree_1198 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2862;
always @( posedge clock ) begin
tree_2862 <= ( $signed( tree_2859 ) ) + ( $signed( tree_2860 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2863;
always @( posedge clock ) begin
tree_2863 <= ( $signed( tree_2861 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2864;
always @( posedge clock ) begin
tree_2864 <= ( $signed( tree_2862 ) ) - ( $signed( tree_2863 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2865;
always @( posedge clock ) begin
tree_2865 <= ( $signed( in[80] ) ) - ( $signed( in[85] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2866;
always @( posedge clock ) begin
tree_2866 <= ( $signed( in[173] ) ) + ( $signed( in[175] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2867;
always @( posedge clock ) begin
tree_2867 <= ( $signed( in[180] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2868;
always @( posedge clock ) begin
tree_2868 <= ( $signed( tree_2865 ) ) - ( $signed( tree_2866 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2869;
always @( posedge clock ) begin
tree_2869 <= ( $signed( tree_2867 ) ) + ( $signed( tree_57 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2870;
always @( posedge clock ) begin
tree_2870 <= ( $signed( tree_89 ) ) + ( $signed( tree_188 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2871;
always @( posedge clock ) begin
tree_2871 <=  - ( $signed( tree_307 ) ) + ( $signed( tree_121 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2872;
always @( posedge clock ) begin
tree_2872 <= ( $signed( tree_308 ) ) - ( $signed( tree_312 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2873;
always @( posedge clock ) begin
tree_2873 <=  - ( $signed( tree_271 ) ) + ( $signed( tree_315 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2874;
always @( posedge clock ) begin
tree_2874 <= ( $signed( tree_325 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2875;
always @( posedge clock ) begin
tree_2875 <= ( $signed( tree_2868 ) ) + ( $signed( tree_2869 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2876;
always @( posedge clock ) begin
tree_2876 <= ( $signed( tree_2870 ) ) + ( $signed( tree_2871 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2877;
always @( posedge clock ) begin
tree_2877 <= ( $signed( tree_2872 ) ) + ( $signed( tree_2873 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2878;
always @( posedge clock ) begin
tree_2878 <= ( $signed( tree_2874 ) ) - ( $signed( tree_310 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2879;
always @( posedge clock ) begin
tree_2879 <= ( $signed( tree_311 ) ) + ( $signed( tree_646 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2880;
always @( posedge clock ) begin
tree_2880 <=  - ( $signed( tree_647 ) ) + ( $signed( tree_314 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2881;
always @( posedge clock ) begin
tree_2881 <= ( $signed( tree_834 ) ) + ( $signed( tree_879 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2882;
always @( posedge clock ) begin
tree_2882 <= ( $signed( tree_318 ) ) + ( $signed( tree_160 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2883;
always @( posedge clock ) begin
tree_2883 <= ( $signed( tree_786 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2884;
always @( posedge clock ) begin
tree_2884 <= ( $signed( tree_2875 ) ) + ( $signed( tree_2876 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2885;
always @( posedge clock ) begin
tree_2885 <= ( $signed( tree_2877 ) ) + ( $signed( tree_2878 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2886;
always @( posedge clock ) begin
tree_2886 <= ( $signed( tree_2879 ) ) + ( $signed( tree_2880 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2887;
always @( posedge clock ) begin
tree_2887 <= ( $signed( tree_2881 ) ) + ( $signed( tree_2882 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2888;
always @( posedge clock ) begin
tree_2888 <=  - ( $signed( tree_2883 ) ) + ( $signed( tree_1108 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2889;
always @( posedge clock ) begin
tree_2889 <= ( $signed( tree_881 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2890;
always @( posedge clock ) begin
tree_2890 <= ( $signed( tree_2884 ) ) + ( $signed( tree_2885 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2891;
always @( posedge clock ) begin
tree_2891 <= ( $signed( tree_2886 ) ) + ( $signed( tree_2887 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2892;
always @( posedge clock ) begin
tree_2892 <= ( $signed( tree_2888 ) ) + ( $signed( tree_2889 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2893;
always @( posedge clock ) begin
tree_2893 <=  - ( $signed( tree_2035 ) ) + ( $signed( tree_886 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2894;
always @( posedge clock ) begin
tree_2894 <= ( $signed( tree_2890 ) ) + ( $signed( tree_2891 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2895;
always @( posedge clock ) begin
tree_2895 <= ( $signed( tree_2892 ) ) + ( $signed( tree_2893 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2896;
always @( posedge clock ) begin
tree_2896 <= ( $signed( tree_2894 ) ) + ( $signed( tree_2895 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2897;
always @( posedge clock ) begin
tree_2897 <= ( $signed( in[70] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2898;
always @( posedge clock ) begin
tree_2898 <=  - ( $signed( tree_2897 ) ) + ( $signed( tree_10 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2899;
always @( posedge clock ) begin
tree_2899 <= ( $signed( tree_39 ) ) + ( $signed( tree_364 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2900;
always @( posedge clock ) begin
tree_2900 <= ( $signed( tree_2898 ) ) - ( $signed( tree_2899 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2901;
always @( posedge clock ) begin
tree_2901 <=  - ( $signed( tree_359 ) ) + ( $signed( tree_361 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2902;
always @( posedge clock ) begin
tree_2902 <= ( $signed( tree_363 ) ) + ( $signed( tree_737 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2903;
always @( posedge clock ) begin
tree_2903 <= ( $signed( tree_911 ) ) - ( $signed( tree_370 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2904;
always @( posedge clock ) begin
tree_2904 <= ( $signed( tree_338 ) ) + ( $signed( tree_372 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2905;
always @( posedge clock ) begin
tree_2905 <= ( $signed( tree_373 ) ) + ( $signed( tree_811 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2906;
always @( posedge clock ) begin
tree_2906 <= ( $signed( tree_914 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2907;
always @( posedge clock ) begin
tree_2907 <= ( $signed( tree_2900 ) ) + ( $signed( tree_2901 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2908;
always @( posedge clock ) begin
tree_2908 <= ( $signed( tree_2902 ) ) + ( $signed( tree_2903 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2909;
always @( posedge clock ) begin
tree_2909 <= ( $signed( tree_2904 ) ) - ( $signed( tree_2905 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2910;
always @( posedge clock ) begin
tree_2910 <=  - ( $signed( tree_2906 ) ) + ( $signed( tree_909 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2911;
always @( posedge clock ) begin
tree_2911 <= ( $signed( tree_368 ) ) + ( $signed( tree_913 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2912;
always @( posedge clock ) begin
tree_2912 <= ( $signed( tree_915 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2913;
always @( posedge clock ) begin
tree_2913 <= ( $signed( tree_2907 ) ) + ( $signed( tree_2908 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2914;
always @( posedge clock ) begin
tree_2914 <= ( $signed( tree_2909 ) ) + ( $signed( tree_2910 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2915;
always @( posedge clock ) begin
tree_2915 <= ( $signed( tree_2911 ) ) + ( $signed( tree_2912 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2916;
always @( posedge clock ) begin
tree_2916 <= ( $signed( tree_2913 ) ) + ( $signed( tree_2914 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2917;
always @( posedge clock ) begin
tree_2917 <= ( $signed( tree_2915 ) ) + ( $signed( tree_2101 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2918;
always @( posedge clock ) begin
tree_2918 <= ( $signed( tree_1209 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2919;
always @( posedge clock ) begin
tree_2919 <= ( $signed( tree_2916 ) ) - ( $signed( tree_2917 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2920;
always @( posedge clock ) begin
tree_2920 <= ( $signed( tree_2918 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2921;
always @( posedge clock ) begin
tree_2921 <= ( $signed( tree_2919 ) ) - ( $signed( tree_2920 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2922;
always @( posedge clock ) begin
tree_2922 <= ( $signed( in[144] ) ) + ( $signed( in[145] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2923;
always @( posedge clock ) begin
tree_2923 <= ( $signed( tree_2922 ) ) + ( $signed( tree_75 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2924;
always @( posedge clock ) begin
tree_2924 <= ( $signed( tree_37 ) ) - ( $signed( tree_26 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2925;
always @( posedge clock ) begin
tree_2925 <= ( $signed( tree_437 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2926;
always @( posedge clock ) begin
tree_2926 <=  - ( $signed( tree_2923 ) ) + ( $signed( tree_2924 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2927;
always @( posedge clock ) begin
tree_2927 <=  - ( $signed( tree_2925 ) ) + ( $signed( tree_45 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2928;
always @( posedge clock ) begin
tree_2928 <= ( $signed( tree_883 ) ) + ( $signed( tree_375 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2929;
always @( posedge clock ) begin
tree_2929 <=  - ( $signed( tree_73 ) ) + ( $signed( tree_310 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2930;
always @( posedge clock ) begin
tree_2930 <= ( $signed( tree_429 ) ) + ( $signed( tree_431 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2931;
always @( posedge clock ) begin
tree_2931 <= ( $signed( tree_2926 ) ) + ( $signed( tree_2927 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2932;
always @( posedge clock ) begin
tree_2932 <= ( $signed( tree_2928 ) ) + ( $signed( tree_2929 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2933;
always @( posedge clock ) begin
tree_2933 <=  - ( $signed( tree_2930 ) ) + ( $signed( tree_428 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2934;
always @( posedge clock ) begin
tree_2934 <= ( $signed( tree_890 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2935;
always @( posedge clock ) begin
tree_2935 <= ( $signed( tree_2931 ) ) + ( $signed( tree_2932 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2936;
always @( posedge clock ) begin
tree_2936 <= ( $signed( tree_2933 ) ) - ( $signed( tree_2934 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2937;
always @( posedge clock ) begin
tree_2937 <= ( $signed( tree_1289 ) ) - ( $signed( tree_1292 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2938;
always @( posedge clock ) begin
tree_2938 <= ( $signed( tree_1293 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2939;
always @( posedge clock ) begin
tree_2939 <= ( $signed( tree_2935 ) ) + ( $signed( tree_2936 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2940;
always @( posedge clock ) begin
tree_2940 <= ( $signed( tree_2937 ) ) - ( $signed( tree_2938 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2941;
always @( posedge clock ) begin
tree_2941 <= ( $signed( tree_2217 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2942;
always @( posedge clock ) begin
tree_2942 <= ( $signed( tree_2939 ) ) + ( $signed( tree_2940 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2943;
always @( posedge clock ) begin
tree_2943 <= ( $signed( tree_2941 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2944;
always @( posedge clock ) begin
tree_2944 <= ( $signed( tree_2942 ) ) + ( $signed( tree_2943 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2945;
always @( posedge clock ) begin
tree_2945 <=  - ( $signed( in[11] ) ) + ( $signed( in[91] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2946;
always @( posedge clock ) begin
tree_2946 <=  - ( $signed( in[124] ) ) + ( $signed( in[125] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2947;
always @( posedge clock ) begin
tree_2947 <= ( $signed( in[136] ) ) - ( $signed( in[158] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2948;
always @( posedge clock ) begin
tree_2948 <= ( $signed( in[191] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2949;
always @( posedge clock ) begin
tree_2949 <= ( $signed( tree_2945 ) ) + ( $signed( tree_2946 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2950;
always @( posedge clock ) begin
tree_2950 <= ( $signed( tree_2947 ) ) - ( $signed( tree_2948 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2951;
always @( posedge clock ) begin
tree_2951 <=  - ( $signed( tree_330 ) ) + ( $signed( tree_489 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2952;
always @( posedge clock ) begin
tree_2952 <=  - ( $signed( tree_351 ) ) + ( $signed( tree_395 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2953;
always @( posedge clock ) begin
tree_2953 <= ( $signed( tree_2949 ) ) + ( $signed( tree_2950 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2954;
always @( posedge clock ) begin
tree_2954 <= ( $signed( tree_2951 ) ) + ( $signed( tree_2952 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2955;
always @( posedge clock ) begin
tree_2955 <= ( $signed( tree_663 ) ) + ( $signed( tree_167 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2956;
always @( posedge clock ) begin
tree_2956 <= ( $signed( tree_1008 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2957;
always @( posedge clock ) begin
tree_2957 <= ( $signed( tree_2953 ) ) + ( $signed( tree_2954 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2958;
always @( posedge clock ) begin
tree_2958 <= ( $signed( tree_2955 ) ) + ( $signed( tree_2956 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2959;
always @( posedge clock ) begin
tree_2959 <= ( $signed( tree_1004 ) ) + ( $signed( tree_1006 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2960;
always @( posedge clock ) begin
tree_2960 <= ( $signed( tree_1212 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2961;
always @( posedge clock ) begin
tree_2961 <= ( $signed( tree_2957 ) ) - ( $signed( tree_2958 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2962;
always @( posedge clock ) begin
tree_2962 <= ( $signed( tree_2959 ) ) + ( $signed( tree_2960 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2963;
always @( posedge clock ) begin
tree_2963 <= ( $signed( tree_1270 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2964;
always @( posedge clock ) begin
tree_2964 <= ( $signed( tree_2961 ) ) + ( $signed( tree_2962 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2965;
always @( posedge clock ) begin
tree_2965 <= ( $signed( tree_2963 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2966;
always @( posedge clock ) begin
tree_2966 <= ( $signed( tree_2964 ) ) - ( $signed( tree_2965 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2967;
always @( posedge clock ) begin
tree_2967 <= ( $signed( tree_2793 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2968;
always @( posedge clock ) begin
tree_2968 <= ( $signed( tree_2966 ) ) - ( $signed( tree_2967 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2969;
always @( posedge clock ) begin
tree_2969 <=  - ( $signed( in[48] ) ) + ( $signed( in[68] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2970;
always @( posedge clock ) begin
tree_2970 <= ( $signed( in[117] ) ) + ( $signed( in[119] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2971;
always @( posedge clock ) begin
tree_2971 <= ( $signed( in[186] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2972;
always @( posedge clock ) begin
tree_2972 <= ( $signed( tree_2969 ) ) + ( $signed( tree_2970 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2973;
always @( posedge clock ) begin
tree_2973 <=  - ( $signed( tree_2971 ) ) + ( $signed( tree_95 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2974;
always @( posedge clock ) begin
tree_2974 <= ( $signed( tree_17 ) ) + ( $signed( tree_264 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2975;
always @( posedge clock ) begin
tree_2975 <= ( $signed( tree_205 ) ) - ( $signed( tree_226 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2976;
always @( posedge clock ) begin
tree_2976 <= ( $signed( tree_2972 ) ) + ( $signed( tree_2973 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2977;
always @( posedge clock ) begin
tree_2977 <=  - ( $signed( tree_2974 ) ) + ( $signed( tree_2975 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2978;
always @( posedge clock ) begin
tree_2978 <= ( $signed( tree_361 ) ) + ( $signed( tree_269 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2979;
always @( posedge clock ) begin
tree_2979 <= ( $signed( tree_257 ) ) - ( $signed( tree_393 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2980;
always @( posedge clock ) begin
tree_2980 <= ( $signed( tree_594 ) ) - ( $signed( tree_596 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2981;
always @( posedge clock ) begin
tree_2981 <= ( $signed( tree_598 ) ) + ( $signed( tree_543 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2982;
always @( posedge clock ) begin
tree_2982 <= ( $signed( tree_472 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2983;
always @( posedge clock ) begin
tree_2983 <= ( $signed( tree_2976 ) ) + ( $signed( tree_2977 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2984;
always @( posedge clock ) begin
tree_2984 <= ( $signed( tree_2978 ) ) + ( $signed( tree_2979 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2985;
always @( posedge clock ) begin
tree_2985 <= ( $signed( tree_2980 ) ) + ( $signed( tree_2981 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2986;
always @( posedge clock ) begin
tree_2986 <= ( $signed( tree_2982 ) ) - ( $signed( tree_1122 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2987;
always @( posedge clock ) begin
tree_2987 <= ( $signed( tree_877 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2988;
always @( posedge clock ) begin
tree_2988 <= ( $signed( tree_2983 ) ) + ( $signed( tree_2984 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2989;
always @( posedge clock ) begin
tree_2989 <= ( $signed( tree_2985 ) ) + ( $signed( tree_2986 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2990;
always @( posedge clock ) begin
tree_2990 <= ( $signed( tree_2987 ) ) + ( $signed( tree_1054 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2991;
always @( posedge clock ) begin
tree_2991 <= ( $signed( tree_977 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2992;
always @( posedge clock ) begin
tree_2992 <= ( $signed( tree_2988 ) ) + ( $signed( tree_2989 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2993;
always @( posedge clock ) begin
tree_2993 <=  - ( $signed( tree_2990 ) ) + ( $signed( tree_2991 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2994;
always @( posedge clock ) begin
tree_2994 <= ( $signed( tree_2465 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2995;
always @( posedge clock ) begin
tree_2995 <= ( $signed( tree_2992 ) ) + ( $signed( tree_2993 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2996;
always @( posedge clock ) begin
tree_2996 <= ( $signed( tree_2994 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2997;
always @( posedge clock ) begin
tree_2997 <= ( $signed( tree_2995 ) ) + ( $signed( tree_2996 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_2998;
always @( posedge clock ) begin
tree_2998 <= ( $signed( in[25] ) ) + ( $signed( in[51] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_2999;
always @( posedge clock ) begin
tree_2999 <= ( $signed( in[125] ) ) + ( $signed( in[148] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3000;
always @( posedge clock ) begin
tree_3000 <= ( $signed( in[156] ) ) + ( $signed( in[173] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3001;
always @( posedge clock ) begin
tree_3001 <= ( $signed( in[188] ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3002;
always @( posedge clock ) begin
tree_3002 <=  - ( $signed( tree_2998 ) ) + ( $signed( tree_2999 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3003;
always @( posedge clock ) begin
tree_3003 <= ( $signed( tree_3000 ) ) + ( $signed( tree_3001 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3004;
always @( posedge clock ) begin
tree_3004 <= ( $signed( tree_21 ) ) + ( $signed( tree_34 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3005;
always @( posedge clock ) begin
tree_3005 <= ( $signed( tree_265 ) ) - ( $signed( tree_97 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3006;
always @( posedge clock ) begin
tree_3006 <=  - ( $signed( tree_632 ) ) + ( $signed( tree_415 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3007;
always @( posedge clock ) begin
tree_3007 <= ( $signed( tree_3002 ) ) + ( $signed( tree_3003 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3008;
always @( posedge clock ) begin
tree_3008 <= ( $signed( tree_3004 ) ) + ( $signed( tree_3005 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3009;
always @( posedge clock ) begin
tree_3009 <= ( $signed( tree_3006 ) ) + ( $signed( tree_645 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3010;
always @( posedge clock ) begin
tree_3010 <=  - ( $signed( tree_641 ) ) + ( $signed( tree_774 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3011;
always @( posedge clock ) begin
tree_3011 <= ( $signed( tree_717 ) ) + ( $signed( tree_705 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_3012;
always @( posedge clock ) begin
tree_3012 <=  - ( $signed( tree_500 ) ) + ( $signed( tree_923 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3013;
always @( posedge clock ) begin
tree_3013 <= ( $signed( tree_3007 ) ) + ( $signed( tree_3008 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3014;
always @( posedge clock ) begin
tree_3014 <= ( $signed( tree_3009 ) ) + ( $signed( tree_3010 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3015;
always @( posedge clock ) begin
tree_3015 <=  - ( $signed( tree_3011 ) ) + ( $signed( tree_3012 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3016;
always @( posedge clock ) begin
tree_3016 <=  - ( $signed( tree_625 ) ) + ( $signed( tree_1151 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3017;
always @( posedge clock ) begin
tree_3017 <= ( $signed( tree_892 ) ) - ( $signed( tree_913 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3018;
always @( posedge clock ) begin
tree_3018 <= ( $signed( tree_3013 ) ) + ( $signed( tree_3014 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3019;
always @( posedge clock ) begin
tree_3019 <= ( $signed( tree_3015 ) ) + ( $signed( tree_3016 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3020;
always @( posedge clock ) begin
tree_3020 <= ( $signed( tree_3017 ) ) - ( $signed( tree_1192 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3021;
always @( posedge clock ) begin
tree_3021 <= ( $signed( tree_980 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_3022;
always @( posedge clock ) begin
tree_3022 <= ( $signed( tree_3018 ) ) + ( $signed( tree_3019 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3023;
always @( posedge clock ) begin
tree_3023 <= ( $signed( tree_3020 ) ) - ( $signed( tree_3021 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3024;
always @( posedge clock ) begin
tree_3024 <= ( $signed( tree_2743 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_3025;
always @( posedge clock ) begin
tree_3025 <= ( $signed( tree_3022 ) ) + ( $signed( tree_3023 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3026;
always @( posedge clock ) begin
tree_3026 <= ( $signed( tree_3024 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_3027;
always @( posedge clock ) begin
tree_3027 <= ( $signed( tree_3025 ) ) - ( $signed( tree_3026 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3028;
always @( posedge clock ) begin
tree_3028 <= ( $signed( in[13] ) ) + ( $signed( in[45] ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_3029;
always @( posedge clock ) begin
tree_3029 <= ( $signed( in[131] ) ) - ( $signed( in[136] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3030;
always @( posedge clock ) begin
tree_3030 <=  - ( $signed( tree_3028 ) ) + ( $signed( tree_3029 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3031;
always @( posedge clock ) begin
tree_3031 <= ( $signed( tree_60 ) ) + ( $signed( tree_61 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_3032;
always @( posedge clock ) begin
tree_3032 <= ( $signed( tree_62 ) ) + ( $signed( tree_66 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3033;
always @( posedge clock ) begin
tree_3033 <= ( $signed( tree_3030 ) ) - ( $signed( tree_3031 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3034;
always @( posedge clock ) begin
tree_3034 <= ( $signed( tree_3032 ) ) + ( $signed( tree_68 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3035;
always @( posedge clock ) begin
tree_3035 <= ( $signed( tree_70 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3036;
always @( posedge clock ) begin
tree_3036 <= ( $signed( tree_3033 ) ) + ( $signed( tree_3034 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3037;
always @( posedge clock ) begin
tree_3037 <= ( $signed( tree_3035 ) ) - ( $signed( tree_1116 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3038;
always @( posedge clock ) begin
tree_3038 <= ( $signed( tree_704 ) ) + ( $signed( tree_1119 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3039;
always @( posedge clock ) begin
tree_3039 <=  - ( $signed( tree_1122 ) ) + ( $signed( tree_710 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3040;
always @( posedge clock ) begin
tree_3040 <= ( $signed( tree_1136 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3041;
always @( posedge clock ) begin
tree_3041 <= ( $signed( tree_3036 ) ) + ( $signed( tree_3037 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3042;
always @( posedge clock ) begin
tree_3042 <= ( $signed( tree_3038 ) ) + ( $signed( tree_3039 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3043;
always @( posedge clock ) begin
tree_3043 <= ( $signed( tree_3040 ) ) + ( $signed( tree_1876 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3044;
always @( posedge clock ) begin
tree_3044 <= ( $signed( tree_1879 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_3045;
always @( posedge clock ) begin
tree_3045 <= ( $signed( tree_3041 ) ) + ( $signed( tree_3042 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3046;
always @( posedge clock ) begin
tree_3046 <= ( $signed( tree_3043 ) ) - ( $signed( tree_3044 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3047;
always @( posedge clock ) begin
tree_3047 <= ( $signed( tree_2742 ) ) + ( $signed( tree_2743 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_3048;
always @( posedge clock ) begin
tree_3048 <= ( $signed( tree_3045 ) ) + ( $signed( tree_3046 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3049;
always @( posedge clock ) begin
tree_3049 <= ( $signed( tree_3047 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_3050;
always @( posedge clock ) begin
tree_3050 <= ( $signed( tree_3048 ) ) - ( $signed( tree_3049 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3051;
always @( posedge clock ) begin
tree_3051 <= ( $signed( in[69] ) ) - ( $signed( in[80] ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3052;
always @( posedge clock ) begin
tree_3052 <= ( $signed( in[154] ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_3053;
always @( posedge clock ) begin
tree_3053 <= ( $signed( tree_3051 ) ) - ( $signed( tree_3052 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3054;
always @( posedge clock ) begin
tree_3054 <= ( $signed( tree_187 ) ) + ( $signed( tree_115 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3055;
always @( posedge clock ) begin
tree_3055 <= ( $signed( tree_1 ) ) + ( $signed( tree_188 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3056;
always @( posedge clock ) begin
tree_3056 <= ( $signed( tree_189 ) ) + ( $signed( tree_190 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_3057;
always @( posedge clock ) begin
tree_3057 <= ( $signed( tree_192 ) ) + ( $signed( tree_193 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3058;
always @( posedge clock ) begin
tree_3058 <= ( $signed( tree_194 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_3059;
always @( posedge clock ) begin
tree_3059 <= ( $signed( tree_3053 ) ) + ( $signed( tree_3054 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3060;
always @( posedge clock ) begin
tree_3060 <= ( $signed( tree_3055 ) ) - ( $signed( tree_3056 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3061;
always @( posedge clock ) begin
tree_3061 <= ( $signed( tree_3057 ) ) - ( $signed( tree_3058 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3062;
always @( posedge clock ) begin
tree_3062 <= ( $signed( tree_86 ) ) - ( $signed( tree_802 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3063;
always @( posedge clock ) begin
tree_3063 <= ( $signed( tree_804 ) ) + ( $signed( tree_806 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_3064;
always @( posedge clock ) begin
tree_3064 <= ( $signed( tree_809 ) ) - ( $signed( tree_811 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3065;
always @( posedge clock ) begin
tree_3065 <= ( $signed( tree_3059 ) ) + ( $signed( tree_3060 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3066;
always @( posedge clock ) begin
tree_3066 <= ( $signed( tree_3061 ) ) + ( $signed( tree_3062 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3067;
always @( posedge clock ) begin
tree_3067 <=  - ( $signed( tree_3063 ) ) + ( $signed( tree_3064 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3068;
always @( posedge clock ) begin
tree_3068 <= ( $signed( tree_1186 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_3069;
always @( posedge clock ) begin
tree_3069 <= ( $signed( tree_3065 ) ) + ( $signed( tree_3066 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3070;
always @( posedge clock ) begin
tree_3070 <= ( $signed( tree_3067 ) ) - ( $signed( tree_3068 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3071;
always @( posedge clock ) begin
tree_3071 <= ( $signed( tree_1182 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3072;
always @( posedge clock ) begin
tree_3072 <= ( $signed( tree_3069 ) ) + ( $signed( tree_3070 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3073;
always @( posedge clock ) begin
tree_3073 <= ( $signed( tree_3071 ) ) - ( $signed( 16'h0 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3074;
always @( posedge clock ) begin
tree_3074 <= ( $signed( tree_3072 ) ) + ( $signed( tree_3073 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] tree_3075;
always @( posedge clock ) begin
tree_3075 <= ( $signed( tree_2793 ) ) + ( $signed( 16'h0 ) ) + ( $signed( 16'h0 ) );
end
reg [15:0] tree_3076;
always @( posedge clock ) begin
tree_3076 <= ( $signed( tree_3074 ) ) - ( $signed( tree_3075 ) ) - ( $signed( 16'h0 ) );
end
reg [15:0] out_0;
assign out[0] = out_0;
reg [15:0] out_1;
assign out[1] = out_1;
assign out[2] = tree_3050;
reg [15:0] out_3;
assign out[3] = out_3;
reg [15:0] out_4;
assign out[4] = out_4;
reg [15:0] out_5;
assign out[5] = out_5;
reg [15:0] out_6;
assign out[6] = out_6;
reg [15:0] out_7;
assign out[7] = out_7;
assign out[8] = tree_3076;
assign out[9] = tree_1997;
assign out[10] = tree_2026;
reg [15:0] out_11;
assign out[11] = out_11;
reg [15:0] out_12;
assign out[12] = out_12;
assign out[13] = tree_2864;
reg [15:0] out_14;
assign out[14] = out_14;
reg [15:0] out_15;
assign out[15] = out_15;
reg [15:0] out_16;
assign out[16] = out_16;
assign out[17] = tree_2096;
assign out[18] = tree_2921;
assign out[19] = tree_2134;
assign out[20] = tree_2164;
reg [15:0] out_21;
assign out[21] = out_21;
reg [15:0] out_22;
assign out[22] = out_22;
assign out[23] = tree_2944;
reg [15:0] out_24;
assign out[24] = out_24;
assign out[25] = tree_2273;
assign out[26] = tree_2309;
reg [15:0] out_27;
assign out[27] = out_27;
reg [15:0] out_28;
assign out[28] = out_28;
assign out[29] = tree_2968;
reg [15:0] out_30;
assign out[30] = out_30;
reg [15:0] out_31;
assign out[31] = out_31;
reg [15:0] out_32;
assign out[32] = out_32;
reg [15:0] out_33;
assign out[33] = out_33;
assign out[34] = tree_2365;
reg [15:0] out_35;
assign out[35] = out_35;
assign out[36] = tree_2396;
assign out[37] = tree_2428;
reg [15:0] out_38;
assign out[38] = out_38;
reg [15:0] out_39;
assign out[39] = out_39;
assign out[40] = tree_2462;
reg [15:0] out_41;
assign out[41] = out_41;
assign out[42] = tree_1584;
assign out[43] = tree_2997;
reg [15:0] out_44;
assign out[44] = out_44;
assign out[45] = tree_2496;
assign out[46] = tree_2524;
assign out[47] = tree_2552;
reg [15:0] out_48;
assign out[48] = out_48;
reg [15:0] out_49;
assign out[49] = out_49;
reg [15:0] out_50;
assign out[50] = out_50;
reg [15:0] out_51;
assign out[51] = out_51;
reg [15:0] out_52;
assign out[52] = out_52;
reg [15:0] out_53;
assign out[53] = out_53;
reg [15:0] out_54;
assign out[54] = out_54;
reg [15:0] out_55;
assign out[55] = out_55;
reg [15:0] out_56;
assign out[56] = out_56;
assign out[57] = tree_2599;
reg [15:0] out_58;
assign out[58] = out_58;
assign out[59] = tree_2631;
reg [15:0] out_60;
assign out[60] = out_60;
reg [15:0] out_61;
assign out[61] = out_61;
assign out[62] = tree_3027;
assign out[63] = tree_2686;
always @( posedge clock ) begin
out_0 <= tree_2712;
out_1 <= tree_2738;
out_3 <= tree_2765;
out_4 <= tree_1905;
out_5 <= tree_2789;
out_6 <= tree_1934;
out_7 <= tree_1961;
out_11 <= tree_2818;
out_12 <= tree_2835;
out_14 <= tree_1257;
out_15 <= tree_2896;
out_16 <= tree_2063;
out_21 <= tree_2190;
out_22 <= tree_2214;
out_24 <= tree_2243;
out_27 <= tree_2334;
out_28 <= tree_1341;
out_30 <= tree_1367;
out_31 <= tree_1392;
out_32 <= tree_1416;
out_33 <= tree_1442;
out_35 <= tree_1472;
out_38 <= tree_1499;
out_39 <= tree_1527;
out_41 <= tree_1557;
out_44 <= tree_1614;
out_48 <= tree_1645;
out_49 <= tree_1674;
out_50 <= tree_1084;
out_51 <= tree_1695;
out_52 <= tree_2574;
out_53 <= tree_1722;
out_54 <= tree_1747;
out_55 <= tree_1775;
out_56 <= tree_1804;
out_58 <= tree_1831;
out_60 <= tree_2652;
out_61 <= tree_1855;
end
endmodule
