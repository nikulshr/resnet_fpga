localparam BN5_CH = 64;
localparam BN5_BW_A = 4;
localparam BN5_BW_B = 15;
localparam BN5_RSHIFT = 8;
localparam BN5_BW_IN = 16;
localparam BN5_BW_OUT = 1;
localparam BN5_MAXVAL = 1;
reg [BN5_CH-1:0][BN5_BW_A-1:0] bn5_a = { 4'h3, 4'h5, 4'h3, 4'h4, 4'h4, 4'h4, 4'h4, 4'h6, 4'h2, 4'h3, 4'h3, 4'h5, 4'h4, 4'h4, 4'h4, 4'h3, 4'h4, 4'h5, 4'h4, 4'h4, 4'h2, 4'h3, 4'h4, 4'h3, 4'h3, 4'h4, 4'h3, 4'h3, 4'h7, 4'h4, 4'h2, 4'h3, 4'h3, 4'h5, 4'h4, 4'h4, 4'h4, 4'h3, 4'h4, 4'h3, 4'h4, 4'h3, 4'h4, 4'h3, 4'h3, 4'h3, 4'h2, 4'h4, 4'h3, 4'h4, 4'h3, 4'h3, 4'h3, 4'h3, 4'h3, 4'h3, 4'h3, 4'h3, 4'h3, 4'h5, 4'h4, 4'h3, 4'h4, 4'h3 };
reg [BN5_CH-1:0][BN5_BW_B-1:0] bn5_b = { 15'h73a9, 15'h722f, 15'h77f1, 15'h7f97, 15'h797a, 15'h75ef, 15'h6822, 15'h6417, 15'h7292, 15'h78c3, 15'h7ee0, 15'h7627, 15'h770e, 15'h026a, 15'h7352, 15'h7561, 15'h7ce6, 15'h754c, 15'h7c50, 15'h4f93, 15'h74c2, 15'h79a6, 15'h7289, 15'h0330, 15'h7752, 15'h0c8c, 15'h7904, 15'h741d, 15'h700d, 15'h6f73, 15'h01f1, 15'h6c6b, 15'h7dbd, 15'h639c, 15'h007d, 15'h7af1, 15'h7cd8, 15'h7c7f, 15'h70b5, 15'h6ac6, 15'h732f, 15'h73ce, 15'h7300, 15'h7fff, 15'h6cf3, 15'h6fad, 15'h7f36, 15'h695f, 15'h6c6b, 15'h761c, 15'h7b70, 15'h74f2, 15'h6bc0, 15'h7b50, 15'h7a31, 15'h06ca, 15'h6d43, 15'h6b33, 15'h7614, 15'h71f7, 15'h6f33, 15'h6852, 15'h08a4, 15'h6a34 };
